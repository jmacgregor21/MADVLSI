magic
tech sky130A
timestamp 1616346938
<< nwell >>
rect 25 920 2120 1620
rect 30 580 2120 920
<< nmos >>
rect 50 0 100 300
rect 150 0 200 300
rect 250 0 300 300
rect 350 0 400 300
rect 450 0 500 300
rect 550 0 600 300
rect 650 0 700 300
rect 750 0 800 300
rect 850 0 900 300
rect 950 0 1000 300
rect 1150 0 1200 300
rect 1250 0 1300 300
rect 1350 0 1400 300
rect 1450 0 1500 300
rect 1550 0 1600 300
rect 1650 0 1700 300
rect 1750 0 1800 300
rect 1850 0 1900 300
rect 1950 0 2000 300
rect 2050 0 2100 300
<< pmos >>
rect 250 1300 300 1600
rect 350 1300 400 1600
rect 450 1300 500 1600
rect 550 1300 600 1600
rect 650 1300 700 1600
rect 750 1300 800 1600
rect 950 1300 1000 1600
rect 1050 1300 1100 1600
rect 1150 1300 1200 1600
rect 1250 1300 1300 1600
rect 1350 1300 1400 1600
rect 1450 1300 1500 1600
rect 1550 1300 1600 1600
rect 1650 1300 1700 1600
rect 1750 1300 1800 1600
rect 1850 1300 1900 1600
rect 150 600 200 900
rect 250 600 300 900
rect 325 600 375 900
rect 425 600 475 900
rect 500 600 550 900
rect 600 600 650 900
rect 675 600 725 900
rect 775 600 825 900
rect 850 600 900 900
rect 950 600 1000 900
rect 1150 600 1200 900
rect 1250 600 1300 900
rect 1325 600 1375 900
rect 1425 600 1475 900
rect 1500 600 1550 900
rect 1600 600 1650 900
rect 1675 600 1725 900
rect 1775 600 1825 900
rect 1850 600 1900 900
rect 1950 600 2000 900
<< ndiff >>
rect 0 285 50 300
rect 0 15 15 285
rect 35 15 50 285
rect 0 0 50 15
rect 100 285 150 300
rect 100 15 115 285
rect 135 15 150 285
rect 100 0 150 15
rect 200 285 250 300
rect 200 15 215 285
rect 235 15 250 285
rect 200 0 250 15
rect 300 285 350 300
rect 300 15 315 285
rect 335 15 350 285
rect 300 0 350 15
rect 400 285 450 300
rect 400 15 415 285
rect 435 15 450 285
rect 400 0 450 15
rect 500 285 550 300
rect 500 15 515 285
rect 535 15 550 285
rect 500 0 550 15
rect 600 285 650 300
rect 600 15 615 285
rect 635 15 650 285
rect 600 0 650 15
rect 700 285 750 300
rect 700 15 715 285
rect 735 15 750 285
rect 700 0 750 15
rect 800 285 850 300
rect 800 15 815 285
rect 835 15 850 285
rect 800 0 850 15
rect 900 285 950 300
rect 900 15 915 285
rect 935 15 950 285
rect 900 0 950 15
rect 1000 285 1050 300
rect 1100 285 1150 300
rect 1000 15 1015 285
rect 1035 15 1050 285
rect 1100 15 1115 285
rect 1135 15 1150 285
rect 1000 0 1050 15
rect 1100 0 1150 15
rect 1200 285 1250 300
rect 1200 15 1215 285
rect 1235 15 1250 285
rect 1200 0 1250 15
rect 1300 285 1350 300
rect 1300 15 1315 285
rect 1335 15 1350 285
rect 1300 0 1350 15
rect 1400 285 1450 300
rect 1400 15 1415 285
rect 1435 15 1450 285
rect 1400 0 1450 15
rect 1500 285 1550 300
rect 1500 15 1515 285
rect 1535 15 1550 285
rect 1500 0 1550 15
rect 1600 285 1650 300
rect 1600 15 1615 285
rect 1635 15 1650 285
rect 1600 0 1650 15
rect 1700 285 1750 300
rect 1700 15 1715 285
rect 1735 15 1750 285
rect 1700 0 1750 15
rect 1800 285 1850 300
rect 1800 15 1815 285
rect 1835 15 1850 285
rect 1800 0 1850 15
rect 1900 285 1950 300
rect 1900 15 1915 285
rect 1935 15 1950 285
rect 1900 0 1950 15
rect 2000 285 2050 300
rect 2000 15 2015 285
rect 2035 15 2050 285
rect 2000 0 2050 15
rect 2100 285 2150 300
rect 2100 15 2115 285
rect 2135 15 2150 285
rect 2100 0 2150 15
<< pdiff >>
rect 200 1585 250 1600
rect 200 1315 215 1585
rect 235 1315 250 1585
rect 200 1300 250 1315
rect 300 1585 350 1600
rect 300 1315 315 1585
rect 335 1315 350 1585
rect 300 1300 350 1315
rect 400 1585 450 1600
rect 400 1315 415 1585
rect 435 1315 450 1585
rect 400 1300 450 1315
rect 500 1585 550 1600
rect 500 1315 515 1585
rect 535 1315 550 1585
rect 500 1300 550 1315
rect 600 1585 650 1600
rect 600 1315 615 1585
rect 635 1315 650 1585
rect 600 1300 650 1315
rect 700 1585 750 1600
rect 700 1315 715 1585
rect 735 1315 750 1585
rect 700 1300 750 1315
rect 800 1585 850 1600
rect 900 1585 950 1600
rect 800 1315 815 1585
rect 835 1315 850 1585
rect 900 1315 915 1585
rect 935 1315 950 1585
rect 800 1300 850 1315
rect 900 1300 950 1315
rect 1000 1585 1050 1600
rect 1000 1315 1015 1585
rect 1035 1315 1050 1585
rect 1000 1300 1050 1315
rect 1100 1585 1150 1600
rect 1100 1315 1115 1585
rect 1135 1315 1150 1585
rect 1100 1300 1150 1315
rect 1200 1585 1250 1600
rect 1200 1315 1215 1585
rect 1235 1315 1250 1585
rect 1200 1300 1250 1315
rect 1300 1585 1350 1600
rect 1300 1315 1315 1585
rect 1335 1315 1350 1585
rect 1300 1300 1350 1315
rect 1400 1585 1450 1600
rect 1400 1315 1415 1585
rect 1435 1315 1450 1585
rect 1400 1300 1450 1315
rect 1500 1585 1550 1600
rect 1500 1315 1515 1585
rect 1535 1315 1550 1585
rect 1500 1300 1550 1315
rect 1600 1585 1650 1600
rect 1600 1315 1615 1585
rect 1635 1315 1650 1585
rect 1600 1300 1650 1315
rect 1700 1585 1750 1600
rect 1700 1315 1715 1585
rect 1735 1315 1750 1585
rect 1700 1300 1750 1315
rect 1800 1585 1850 1600
rect 1800 1315 1815 1585
rect 1835 1315 1850 1585
rect 1800 1300 1850 1315
rect 1900 1585 1950 1600
rect 1900 1315 1915 1585
rect 1935 1315 1950 1585
rect 1900 1300 1950 1315
rect 100 885 150 900
rect 100 615 115 885
rect 135 615 150 885
rect 100 600 150 615
rect 200 885 250 900
rect 200 615 215 885
rect 235 615 250 885
rect 200 600 250 615
rect 300 600 325 900
rect 375 885 425 900
rect 375 615 390 885
rect 410 615 425 885
rect 375 600 425 615
rect 475 600 500 900
rect 550 885 600 900
rect 550 615 565 885
rect 585 615 600 885
rect 550 600 600 615
rect 650 600 675 900
rect 725 885 775 900
rect 725 615 740 885
rect 760 615 775 885
rect 725 600 775 615
rect 825 600 850 900
rect 900 885 950 900
rect 900 615 915 885
rect 935 615 950 885
rect 900 600 950 615
rect 1000 885 1050 900
rect 1100 885 1150 900
rect 1000 615 1015 885
rect 1035 615 1050 885
rect 1100 615 1115 885
rect 1135 615 1150 885
rect 1000 600 1050 615
rect 1100 600 1150 615
rect 1200 885 1250 900
rect 1200 615 1215 885
rect 1235 615 1250 885
rect 1200 600 1250 615
rect 1300 600 1325 900
rect 1375 885 1425 900
rect 1375 615 1390 885
rect 1410 615 1425 885
rect 1375 600 1425 615
rect 1475 600 1500 900
rect 1550 885 1600 900
rect 1550 615 1565 885
rect 1585 615 1600 885
rect 1550 600 1600 615
rect 1650 600 1675 900
rect 1725 885 1775 900
rect 1725 615 1740 885
rect 1760 615 1775 885
rect 1725 600 1775 615
rect 1825 600 1850 900
rect 1900 885 1950 900
rect 1900 615 1915 885
rect 1935 615 1950 885
rect 1900 600 1950 615
rect 2000 885 2050 900
rect 2000 615 2015 885
rect 2035 615 2050 885
rect 2000 600 2050 615
<< ndiffc >>
rect 15 15 35 285
rect 115 15 135 285
rect 215 15 235 285
rect 315 15 335 285
rect 415 15 435 285
rect 515 15 535 285
rect 615 15 635 285
rect 715 15 735 285
rect 815 15 835 285
rect 915 15 935 285
rect 1015 15 1035 285
rect 1115 15 1135 285
rect 1215 15 1235 285
rect 1315 15 1335 285
rect 1415 15 1435 285
rect 1515 15 1535 285
rect 1615 15 1635 285
rect 1715 15 1735 285
rect 1815 15 1835 285
rect 1915 15 1935 285
rect 2015 15 2035 285
rect 2115 15 2135 285
<< pdiffc >>
rect 215 1315 235 1585
rect 315 1315 335 1585
rect 415 1315 435 1585
rect 515 1315 535 1585
rect 615 1315 635 1585
rect 715 1315 735 1585
rect 815 1315 835 1585
rect 915 1315 935 1585
rect 1015 1315 1035 1585
rect 1115 1315 1135 1585
rect 1215 1315 1235 1585
rect 1315 1315 1335 1585
rect 1415 1315 1435 1585
rect 1515 1315 1535 1585
rect 1615 1315 1635 1585
rect 1715 1315 1735 1585
rect 1815 1315 1835 1585
rect 1915 1315 1935 1585
rect 115 615 135 885
rect 215 615 235 885
rect 390 615 410 885
rect 565 615 585 885
rect 740 615 760 885
rect 915 615 935 885
rect 1015 615 1035 885
rect 1115 615 1135 885
rect 1215 615 1235 885
rect 1390 615 1410 885
rect 1565 615 1585 885
rect 1740 615 1760 885
rect 1915 615 1935 885
rect 2015 615 2035 885
<< psubdiff >>
rect -50 285 0 300
rect -50 15 -35 285
rect -15 15 0 285
rect -50 0 0 15
rect 1050 285 1100 300
rect 1050 15 1065 285
rect 1085 15 1100 285
rect 1050 0 1100 15
rect 2150 285 2200 300
rect 2150 15 2165 285
rect 2185 15 2200 285
rect 2150 0 2200 15
<< nsubdiff >>
rect 150 1585 200 1600
rect 150 1315 165 1585
rect 185 1315 200 1585
rect 150 1300 200 1315
rect 850 1585 900 1600
rect 850 1315 865 1585
rect 885 1315 900 1585
rect 850 1300 900 1315
rect 1950 1585 2000 1600
rect 1950 1315 1965 1585
rect 1985 1315 2000 1585
rect 1950 1300 2000 1315
rect 50 885 100 900
rect 50 615 65 885
rect 85 615 100 885
rect 50 600 100 615
rect 1050 885 1100 900
rect 1050 615 1065 885
rect 1085 615 1100 885
rect 1050 600 1100 615
rect 2050 885 2100 900
rect 2050 615 2065 885
rect 2085 615 2100 885
rect 2050 600 2100 615
<< psubdiffcont >>
rect -35 15 -15 285
rect 1065 15 1085 285
rect 2165 15 2185 285
<< nsubdiffcont >>
rect 165 1315 185 1585
rect 865 1315 885 1585
rect 1965 1315 1985 1585
rect 65 615 85 885
rect 1065 615 1085 885
rect 2065 615 2085 885
<< poly >>
rect 25 1745 1200 1760
rect 1150 1730 1700 1745
rect 25 1705 1100 1720
rect 1050 1690 1100 1705
rect 245 1670 285 1680
rect 245 1650 255 1670
rect 275 1650 285 1670
rect 245 1640 285 1650
rect 1050 1670 1065 1690
rect 1085 1670 1100 1690
rect 250 1615 265 1640
rect 250 1600 300 1615
rect 350 1600 400 1615
rect 450 1600 500 1615
rect 550 1600 600 1615
rect 650 1600 700 1615
rect 750 1600 800 1615
rect 950 1600 1000 1640
rect 1050 1600 1100 1670
rect 1150 1600 1200 1730
rect 1250 1600 1300 1730
rect 1350 1690 1400 1705
rect 1350 1670 1365 1690
rect 1385 1670 1400 1690
rect 1350 1600 1400 1670
rect 1450 1690 1500 1705
rect 1450 1670 1465 1690
rect 1485 1670 1500 1690
rect 1450 1600 1500 1670
rect 1550 1600 1600 1730
rect 1650 1600 1700 1730
rect 1750 1690 1800 1705
rect 1750 1670 1765 1690
rect 1785 1670 1800 1690
rect 1750 1600 1800 1670
rect 1860 1650 1900 1660
rect 1860 1630 1870 1650
rect 1890 1630 1900 1650
rect 1860 1615 1900 1630
rect 1850 1600 1900 1615
rect 250 1285 300 1300
rect 350 1285 400 1300
rect 450 1285 500 1300
rect 550 1285 600 1300
rect 650 1285 700 1300
rect 350 1270 700 1285
rect 750 1285 800 1300
rect 950 1285 1000 1300
rect 1050 1285 1100 1300
rect 1150 1285 1200 1300
rect 1250 1285 1300 1300
rect 1350 1285 1400 1300
rect 1450 1285 1500 1300
rect 1550 1285 1600 1300
rect 1650 1285 1700 1300
rect 1750 1285 1800 1300
rect 1850 1285 1900 1300
rect 750 1275 1000 1285
rect 750 1270 865 1275
rect 350 1260 395 1270
rect 25 1245 395 1260
rect 855 1255 865 1270
rect 885 1270 1000 1275
rect 885 1255 895 1270
rect 855 1245 895 1255
rect 1205 1250 1245 1260
rect 1205 1230 1215 1250
rect 1235 1235 1245 1250
rect 1605 1250 1645 1260
rect 1605 1235 1615 1250
rect 1235 1230 1615 1235
rect 1635 1235 1645 1250
rect 1635 1230 2135 1235
rect 1205 1220 2135 1230
rect 0 1000 1825 1015
rect 250 965 300 975
rect 150 945 190 955
rect 150 925 160 945
rect 180 925 190 945
rect 150 915 190 925
rect 250 945 265 965
rect 285 945 300 965
rect 150 900 200 915
rect 250 900 300 945
rect 325 900 375 1000
rect 425 900 475 1000
rect 500 965 550 975
rect 500 945 515 965
rect 535 945 550 965
rect 500 900 550 945
rect 600 965 650 975
rect 600 945 615 965
rect 635 945 650 965
rect 600 900 650 945
rect 675 900 725 1000
rect 775 900 825 1000
rect 850 965 900 975
rect 850 945 865 965
rect 885 945 900 965
rect 850 900 900 945
rect 1250 955 1300 970
rect 1250 935 1265 955
rect 1285 935 1300 955
rect 950 900 1000 915
rect 1150 900 1200 915
rect 1250 900 1300 935
rect 1325 900 1375 1000
rect 1425 900 1475 1000
rect 1500 955 1550 970
rect 1500 935 1515 955
rect 1535 935 1550 955
rect 1500 900 1550 935
rect 1600 955 1650 970
rect 1600 935 1615 955
rect 1635 935 1650 955
rect 1600 900 1650 935
rect 1675 900 1725 1000
rect 1775 900 1825 1000
rect 1850 955 1900 970
rect 1850 935 1865 955
rect 1885 935 1900 955
rect 1850 900 1900 935
rect 1950 955 2000 970
rect 1950 935 1965 955
rect 1985 935 2000 955
rect 1950 900 2000 935
rect 150 585 200 600
rect 250 585 300 600
rect 325 585 375 600
rect 425 585 475 600
rect 500 585 550 600
rect 600 585 650 600
rect 675 585 725 600
rect 775 585 825 600
rect 850 585 900 600
rect 950 585 1000 600
rect 1055 585 1095 590
rect 1150 585 1200 600
rect 1250 585 1300 600
rect 1325 585 1375 600
rect 1425 585 1475 600
rect 1500 585 1550 600
rect 1600 585 1650 600
rect 1675 585 1725 600
rect 1775 585 1825 600
rect 1850 585 1900 600
rect 1950 585 2000 600
rect 950 580 1200 585
rect 950 570 1065 580
rect 1055 560 1065 570
rect 1085 570 1200 580
rect 1085 560 1095 570
rect 1055 550 1095 560
rect -70 510 265 525
rect 130 475 170 485
rect 130 455 140 475
rect 160 455 170 475
rect 130 445 170 455
rect 130 380 145 445
rect 105 370 145 380
rect 5 345 45 355
rect 5 325 15 345
rect 35 330 45 345
rect 105 350 115 370
rect 135 350 145 370
rect 105 340 145 350
rect 250 395 265 510
rect 2120 460 2135 1220
rect 1905 450 2135 460
rect 1905 430 1915 450
rect 1935 445 2135 450
rect 1935 430 1945 445
rect 1905 420 1945 430
rect 250 380 1900 395
rect 35 325 70 330
rect 5 315 70 325
rect 50 300 100 315
rect 150 300 200 315
rect 250 300 300 380
rect 350 300 400 380
rect 450 300 500 315
rect 550 300 600 315
rect 650 300 700 380
rect 750 300 800 380
rect 1055 345 1095 355
rect 1055 330 1065 345
rect 950 325 1065 330
rect 1085 330 1095 345
rect 1085 325 1200 330
rect 950 315 1200 325
rect 850 300 900 315
rect 950 300 1000 315
rect 1150 300 1200 315
rect 1250 300 1300 315
rect 1350 300 1400 380
rect 1450 300 1500 380
rect 1550 300 1600 315
rect 1650 300 1700 315
rect 1750 300 1800 380
rect 1850 300 1900 380
rect 2060 355 2100 365
rect 2060 335 2070 355
rect 2090 335 2100 355
rect 2060 315 2100 335
rect 1950 300 2000 315
rect 2050 300 2100 315
rect 50 -15 100 0
rect 150 -40 200 0
rect 250 -15 300 0
rect 350 -15 400 0
rect 450 -40 500 0
rect 550 -40 600 0
rect 650 -15 700 0
rect 750 -15 800 0
rect 850 -40 900 0
rect 950 -15 1000 0
rect 1150 -15 1200 0
rect 1250 -40 1300 0
rect 1350 -15 1400 0
rect 1450 -15 1500 0
rect 1550 -40 1600 0
rect 1650 -40 1700 0
rect 1750 -15 1800 0
rect 1850 -15 1900 0
rect 1950 -40 2000 0
rect 2050 -15 2100 0
rect -70 -55 2000 -40
<< polycont >>
rect 255 1650 275 1670
rect 1065 1670 1085 1690
rect 1365 1670 1385 1690
rect 1465 1670 1485 1690
rect 1765 1670 1785 1690
rect 1870 1630 1890 1650
rect 865 1255 885 1275
rect 1215 1230 1235 1250
rect 1615 1230 1635 1250
rect 160 925 180 945
rect 265 945 285 965
rect 515 945 535 965
rect 615 945 635 965
rect 865 945 885 965
rect 1265 935 1285 955
rect 1515 935 1535 955
rect 1615 935 1635 955
rect 1865 935 1885 955
rect 1965 935 1985 955
rect 1065 560 1085 580
rect 140 455 160 475
rect 15 325 35 345
rect 115 350 135 370
rect 1915 430 1935 450
rect 1065 325 1085 345
rect 2070 335 2090 355
<< locali >>
rect 1055 1690 1795 1700
rect 245 1670 285 1680
rect 245 1660 255 1670
rect 225 1650 255 1660
rect 275 1650 285 1670
rect 1055 1670 1065 1690
rect 1085 1670 1365 1690
rect 1385 1670 1465 1690
rect 1485 1670 1765 1690
rect 1785 1670 1795 1690
rect 1055 1660 1795 1670
rect 225 1640 285 1650
rect 1860 1650 1900 1660
rect 225 1595 245 1640
rect 155 1585 245 1595
rect 155 1315 165 1585
rect 185 1315 215 1585
rect 235 1315 245 1585
rect 155 1305 245 1315
rect 305 1620 1745 1640
rect 1860 1630 1870 1650
rect 1890 1640 1900 1650
rect 1890 1630 1925 1640
rect 1860 1620 1925 1630
rect 305 1585 345 1620
rect 305 1315 315 1585
rect 335 1315 345 1585
rect 305 1305 345 1315
rect 405 1585 445 1595
rect 405 1315 415 1585
rect 435 1315 445 1585
rect 405 1305 445 1315
rect 505 1585 545 1620
rect 505 1315 515 1585
rect 535 1315 545 1585
rect 505 1305 545 1315
rect 605 1585 645 1595
rect 605 1315 615 1585
rect 635 1315 645 1585
rect 605 1305 645 1315
rect 705 1585 745 1620
rect 705 1315 715 1585
rect 735 1315 745 1585
rect 705 1305 745 1315
rect 805 1585 945 1595
rect 805 1315 815 1585
rect 835 1315 865 1585
rect 885 1315 915 1585
rect 935 1315 945 1585
rect 805 1305 945 1315
rect 1005 1585 1045 1595
rect 1005 1315 1015 1585
rect 1035 1315 1045 1585
rect 855 1275 895 1305
rect 855 1255 865 1275
rect 885 1255 895 1275
rect 855 1245 895 1255
rect 1005 1200 1045 1315
rect 1105 1585 1145 1620
rect 1105 1315 1115 1585
rect 1135 1315 1145 1585
rect 1105 1305 1145 1315
rect 1205 1585 1245 1595
rect 1205 1315 1215 1585
rect 1235 1315 1245 1585
rect 1205 1250 1245 1315
rect 1305 1585 1345 1620
rect 1305 1315 1315 1585
rect 1335 1315 1345 1585
rect 1305 1305 1345 1315
rect 1405 1585 1445 1595
rect 1405 1315 1415 1585
rect 1435 1315 1445 1585
rect 1205 1230 1215 1250
rect 1235 1230 1245 1250
rect 1205 1220 1245 1230
rect 1405 1200 1445 1315
rect 1505 1585 1545 1620
rect 1505 1315 1515 1585
rect 1535 1315 1545 1585
rect 1505 1305 1545 1315
rect 1605 1585 1645 1595
rect 1605 1315 1615 1585
rect 1635 1315 1645 1585
rect 1605 1250 1645 1315
rect 1705 1585 1745 1620
rect 1905 1595 1925 1620
rect 1705 1315 1715 1585
rect 1735 1315 1745 1585
rect 1705 1305 1745 1315
rect 1805 1585 1845 1595
rect 1805 1315 1815 1585
rect 1835 1315 1845 1585
rect 1605 1230 1615 1250
rect 1635 1230 1645 1250
rect 1605 1220 1645 1230
rect 1805 1200 1845 1315
rect 1905 1585 1995 1595
rect 1905 1315 1915 1585
rect 1935 1315 1965 1585
rect 1985 1315 1995 1585
rect 1905 1305 1995 1315
rect 5 1180 1845 1200
rect 5 425 25 1180
rect 255 965 900 975
rect 150 945 190 955
rect 150 935 160 945
rect 125 925 160 935
rect 180 925 190 945
rect 255 945 265 965
rect 285 945 515 965
rect 535 945 615 965
rect 635 945 865 965
rect 885 960 900 965
rect 1255 960 1895 965
rect 885 955 1895 960
rect 885 945 1265 955
rect 255 935 1265 945
rect 1285 935 1515 955
rect 1535 935 1615 955
rect 1635 935 1865 955
rect 1885 935 1895 955
rect 125 915 190 925
rect 125 895 145 915
rect 55 885 145 895
rect 55 615 65 885
rect 85 615 115 885
rect 135 615 145 885
rect 55 605 145 615
rect 205 885 245 895
rect 205 615 215 885
rect 235 615 245 885
rect 205 605 245 615
rect 380 885 420 935
rect 380 615 390 885
rect 410 615 420 885
rect 380 560 420 615
rect 555 885 595 895
rect 555 615 565 885
rect 585 615 595 885
rect 555 605 595 615
rect 730 885 770 935
rect 1255 925 1895 935
rect 1955 955 2025 965
rect 1955 935 1965 955
rect 1985 935 2025 955
rect 1955 925 2025 935
rect 2005 895 2025 925
rect 730 615 740 885
rect 760 615 770 885
rect 730 560 770 615
rect 905 885 945 895
rect 905 615 915 885
rect 935 615 945 885
rect 905 605 945 615
rect 1005 885 1145 895
rect 1005 615 1015 885
rect 1035 615 1065 885
rect 1085 615 1115 885
rect 1135 615 1145 885
rect 1005 605 1145 615
rect 1205 885 1245 895
rect 1205 615 1215 885
rect 1235 615 1245 885
rect 1205 605 1245 615
rect 1380 885 1420 895
rect 1380 615 1390 885
rect 1410 615 1420 885
rect 150 540 770 560
rect 1055 580 1095 605
rect 1055 560 1065 580
rect 1085 560 1095 580
rect 1380 580 1420 615
rect 1555 885 1595 895
rect 1555 615 1565 885
rect 1585 615 1595 885
rect 1555 605 1595 615
rect 1730 885 1770 895
rect 1730 615 1740 885
rect 1760 615 1770 885
rect 1730 580 1770 615
rect 1905 885 1945 895
rect 1905 615 1915 885
rect 1935 615 1945 885
rect 1905 605 1945 615
rect 2005 885 2095 895
rect 2005 615 2015 885
rect 2035 615 2065 885
rect 2085 615 2095 885
rect 2005 605 2095 615
rect 1380 560 2025 580
rect 1055 550 1095 560
rect 150 485 170 540
rect 130 475 170 485
rect 130 455 140 475
rect 160 455 170 475
rect 2005 460 2025 560
rect 130 445 170 455
rect 1905 450 1945 460
rect 1905 430 1915 450
rect 1935 430 1945 450
rect 5 405 245 425
rect 105 370 145 380
rect 5 345 45 355
rect 5 325 15 345
rect 35 325 45 345
rect 5 315 45 325
rect 25 295 45 315
rect -45 285 45 295
rect -45 15 -35 285
rect -15 15 15 285
rect 35 15 45 285
rect -45 5 45 15
rect 105 350 115 370
rect 135 350 145 370
rect 105 285 145 350
rect 105 15 115 285
rect 135 15 145 285
rect 105 -20 145 15
rect 205 340 245 405
rect 1055 345 1095 355
rect 205 320 845 340
rect 205 285 245 320
rect 205 15 215 285
rect 235 15 245 285
rect 205 5 245 15
rect 305 285 345 295
rect 305 15 315 285
rect 335 15 345 285
rect 305 5 345 15
rect 405 285 445 320
rect 405 15 415 285
rect 435 15 445 285
rect 405 5 445 15
rect 505 285 545 295
rect 505 15 515 285
rect 535 15 545 285
rect 505 -20 545 15
rect 605 285 645 320
rect 605 15 615 285
rect 635 15 645 285
rect 605 5 645 15
rect 705 285 745 295
rect 705 15 715 285
rect 735 15 745 285
rect 705 5 745 15
rect 805 285 845 320
rect 1055 325 1065 345
rect 1085 325 1095 345
rect 1905 340 1945 430
rect 1055 295 1095 325
rect 1305 320 1945 340
rect 805 15 815 285
rect 835 15 845 285
rect 805 5 845 15
rect 905 285 945 295
rect 905 15 915 285
rect 935 15 945 285
rect 905 -20 945 15
rect 1005 285 1145 295
rect 1005 15 1015 285
rect 1035 15 1065 285
rect 1085 15 1115 285
rect 1135 15 1145 285
rect 1005 5 1145 15
rect 1205 285 1245 295
rect 1205 15 1215 285
rect 1235 15 1245 285
rect 105 -40 945 -20
rect 1205 -15 1245 15
rect 1305 285 1345 320
rect 1305 15 1315 285
rect 1335 15 1345 285
rect 1305 5 1345 15
rect 1405 285 1445 295
rect 1405 15 1415 285
rect 1435 15 1445 285
rect 1405 5 1445 15
rect 1505 285 1545 320
rect 1505 15 1515 285
rect 1535 15 1545 285
rect 1505 5 1545 15
rect 1605 285 1645 295
rect 1605 15 1615 285
rect 1635 15 1645 285
rect 1605 -15 1645 15
rect 1705 285 1745 320
rect 1705 15 1715 285
rect 1735 15 1745 285
rect 1705 5 1745 15
rect 1805 285 1845 295
rect 1805 15 1815 285
rect 1835 15 1845 285
rect 1805 5 1845 15
rect 1905 285 1945 320
rect 1905 15 1915 285
rect 1935 15 1945 285
rect 1905 5 1945 15
rect 2005 440 2220 460
rect 2005 315 2025 440
rect 2060 355 2145 365
rect 2060 335 2070 355
rect 2090 335 2145 355
rect 2060 325 2145 335
rect 2005 285 2045 315
rect 2005 15 2015 285
rect 2035 15 2045 285
rect 2005 -15 2045 15
rect 2105 295 2145 325
rect 2105 285 2195 295
rect 2105 15 2115 285
rect 2135 15 2165 285
rect 2185 15 2195 285
rect 2105 5 2195 15
rect 1205 -35 2045 -15
<< viali >>
rect 165 1315 185 1585
rect 215 1315 235 1585
rect 415 1315 435 1585
rect 615 1315 635 1585
rect 815 1315 835 1585
rect 865 1315 885 1585
rect 915 1315 935 1585
rect 1915 1315 1935 1585
rect 1965 1315 1985 1585
rect 65 615 85 885
rect 115 615 135 885
rect 215 615 235 885
rect 565 615 585 885
rect 915 615 935 885
rect 1015 615 1035 885
rect 1065 615 1085 885
rect 1115 615 1135 885
rect 1215 615 1235 885
rect 1565 615 1585 885
rect 1915 615 1935 885
rect 2015 615 2035 885
rect 2065 615 2085 885
rect -35 15 -15 285
rect 15 15 35 285
rect 315 15 335 285
rect 715 15 735 285
rect 1015 15 1035 285
rect 1065 15 1085 285
rect 1115 15 1135 285
rect 1415 15 1435 285
rect 1815 15 1835 285
rect 2115 15 2135 285
rect 2165 15 2185 285
<< metal1 >>
rect 25 1585 2120 1605
rect 25 1315 165 1585
rect 185 1315 215 1585
rect 235 1315 415 1585
rect 435 1315 615 1585
rect 635 1315 815 1585
rect 835 1315 865 1585
rect 885 1315 915 1585
rect 935 1315 1915 1585
rect 1935 1315 1965 1585
rect 1985 1315 2120 1585
rect 25 885 2120 1315
rect 25 615 65 885
rect 85 615 115 885
rect 135 615 215 885
rect 235 615 565 885
rect 585 615 915 885
rect 935 615 1015 885
rect 1035 615 1065 885
rect 1085 615 1115 885
rect 1135 615 1215 885
rect 1235 615 1565 885
rect 1585 615 1915 885
rect 1935 615 2015 885
rect 2035 615 2065 885
rect 2085 615 2120 885
rect 25 600 2120 615
rect -70 285 2220 300
rect -70 15 -35 285
rect -15 15 15 285
rect 35 15 315 285
rect 335 15 715 285
rect 735 15 1015 285
rect 1035 15 1065 285
rect 1085 15 1115 285
rect 1135 15 1415 285
rect 1435 15 1815 285
rect 1835 15 2115 285
rect 2135 15 2165 285
rect 2185 15 2220 285
rect -70 0 2220 15
<< labels >>
rlabel poly 25 1750 25 1750 7 V2
port 2 w
rlabel poly 25 1710 25 1710 7 V1
port 1 w
rlabel locali 2220 450 2220 450 3 Vout
port 9 e
rlabel poly -70 515 -70 515 7 Vbn
port 8 w
rlabel poly -70 -50 -70 -50 7 Vcn
port 7 w
rlabel poly 25 1250 25 1250 7 Vbp
port 6 w
rlabel poly 0 1005 0 1005 7 Vcp
port 5 w
rlabel metal1 25 1485 25 1485 7 VP
port 3 w
rlabel pdiff 1830 700 1830 700 7 net12
rlabel pdiff 1665 705 1665 705 7 net11
rlabel pdiff 310 690 310 690 7 net4
rlabel pdiff 490 685 490 685 7 net5
rlabel pdiff 660 680 660 680 7 net6
rlabel metal1 -70 205 -70 205 7 VN
port 4 w
rlabel locali 440 545 440 545 7 net8
<< end >>
