magic
tech sky130A
timestamp 1616270437
<< nwell >>
rect -120 1480 3195 1820
rect -320 980 3470 1320
<< nmos >>
rect 0 500 50 800
rect 100 500 150 800
rect 200 500 250 800
rect 300 500 350 800
rect 400 500 450 800
rect 500 500 550 800
rect 600 500 650 800
rect 700 500 750 800
rect 800 500 850 800
rect 900 500 950 800
rect 1000 500 1050 800
rect 1100 500 1150 800
rect 1200 500 1250 800
rect 1300 500 1350 800
rect 1400 500 1450 800
rect 1500 500 1550 800
rect 1600 500 1650 800
rect 1700 500 1750 800
rect 1800 500 1850 800
rect 1900 500 1950 800
rect 2000 500 2050 800
rect 2100 500 2150 800
rect 2300 500 2350 800
rect 2400 500 2450 800
rect 2500 500 2550 800
rect 2600 500 2650 800
rect 2700 500 2750 800
rect 2800 500 2850 800
rect 0 0 50 300
rect 100 0 150 300
rect 200 0 250 300
rect 300 0 350 300
rect 400 0 450 300
rect 500 0 550 300
rect 700 0 750 300
rect 800 0 850 300
rect 875 0 925 300
rect 950 0 1000 300
rect 1025 0 1075 300
rect 1100 0 1150 300
rect 1175 0 1225 300
rect 1250 0 1300 300
rect 1325 0 1375 300
rect 1400 0 1450 300
rect 1475 0 1525 300
rect 1550 0 1600 300
rect 1625 0 1675 300
rect 1700 0 1750 300
rect 1775 0 1825 300
rect 1850 0 1900 300
rect 1925 0 1975 300
rect 2000 0 2050 300
rect 2075 0 2125 300
rect 2150 0 2200 300
rect 2225 0 2275 300
rect 2325 0 2375 300
rect 2525 0 2575 300
rect 2625 0 2675 300
rect 2725 0 2775 300
rect 2825 0 2875 300
rect 2925 0 2975 300
rect 3025 0 3075 300
<< pmos >>
rect 0 1500 50 1800
rect 100 1500 150 1800
rect 200 1500 250 1800
rect 300 1500 350 1800
rect 400 1500 450 1800
rect 500 1500 550 1800
rect 700 1500 750 1800
rect 800 1500 850 1800
rect 875 1500 925 1800
rect 950 1500 1000 1800
rect 1025 1500 1075 1800
rect 1100 1500 1150 1800
rect 1175 1500 1225 1800
rect 1250 1500 1300 1800
rect 1325 1500 1375 1800
rect 1400 1500 1450 1800
rect 1475 1500 1525 1800
rect 1550 1500 1600 1800
rect 1625 1500 1675 1800
rect 1700 1500 1750 1800
rect 1775 1500 1825 1800
rect 1850 1500 1900 1800
rect 1925 1500 1975 1800
rect 2000 1500 2050 1800
rect 2075 1500 2125 1800
rect 2150 1500 2200 1800
rect 2225 1500 2275 1800
rect 2325 1500 2375 1800
rect 2525 1500 2575 1800
rect 2625 1500 2675 1800
rect 2725 1500 2775 1800
rect 2825 1500 2875 1800
rect 2925 1500 2975 1800
rect 3025 1500 3075 1800
rect -200 1000 -150 1300
rect -100 1000 -50 1300
rect 0 1000 50 1300
rect 100 1000 150 1300
rect 200 1000 250 1300
rect 300 1000 350 1300
rect 500 1000 550 1300
rect 600 1000 650 1300
rect 700 1000 750 1300
rect 800 1000 850 1300
rect 900 1000 950 1300
rect 1000 1000 1050 1300
rect 1100 1000 1150 1300
rect 1200 1000 1250 1300
rect 1300 1000 1350 1300
rect 1400 1000 1450 1300
rect 1500 1000 1550 1300
rect 1600 1000 1650 1300
rect 1700 1000 1750 1300
rect 1800 1000 1850 1300
rect 1900 1000 1950 1300
rect 2000 1000 2050 1300
rect 2100 1000 2150 1300
rect 2200 1000 2250 1300
rect 2300 1000 2350 1300
rect 2400 1000 2450 1300
rect 2500 1000 2550 1300
rect 2600 1000 2650 1300
rect 2800 1000 2850 1300
rect 2900 1000 2950 1300
rect 3000 1000 3050 1300
rect 3100 1000 3150 1300
rect 3200 1000 3250 1300
rect 3300 1000 3350 1300
<< ndiff >>
rect -50 785 0 800
rect -50 515 -35 785
rect -15 515 0 785
rect -50 500 0 515
rect 50 785 100 800
rect 50 515 65 785
rect 85 515 100 785
rect 50 500 100 515
rect 150 785 200 800
rect 150 515 165 785
rect 185 515 200 785
rect 150 500 200 515
rect 250 785 300 800
rect 250 515 265 785
rect 285 515 300 785
rect 250 500 300 515
rect 350 785 400 800
rect 350 515 365 785
rect 385 515 400 785
rect 350 500 400 515
rect 450 785 500 800
rect 450 515 465 785
rect 485 515 500 785
rect 450 500 500 515
rect 550 785 600 800
rect 550 515 565 785
rect 585 515 600 785
rect 550 500 600 515
rect 650 785 700 800
rect 650 515 665 785
rect 685 515 700 785
rect 650 500 700 515
rect 750 785 800 800
rect 750 515 765 785
rect 785 515 800 785
rect 750 500 800 515
rect 850 785 900 800
rect 850 515 865 785
rect 885 515 900 785
rect 850 500 900 515
rect 950 785 1000 800
rect 950 515 965 785
rect 985 515 1000 785
rect 950 500 1000 515
rect 1050 785 1100 800
rect 1050 515 1065 785
rect 1085 515 1100 785
rect 1050 500 1100 515
rect 1150 785 1200 800
rect 1150 515 1165 785
rect 1185 515 1200 785
rect 1150 500 1200 515
rect 1250 785 1300 800
rect 1250 515 1265 785
rect 1285 515 1300 785
rect 1250 500 1300 515
rect 1350 785 1400 800
rect 1350 515 1365 785
rect 1385 515 1400 785
rect 1350 500 1400 515
rect 1450 785 1500 800
rect 1450 515 1465 785
rect 1485 515 1500 785
rect 1450 500 1500 515
rect 1550 785 1600 800
rect 1550 515 1565 785
rect 1585 515 1600 785
rect 1550 500 1600 515
rect 1650 785 1700 800
rect 1650 515 1665 785
rect 1685 515 1700 785
rect 1650 500 1700 515
rect 1750 785 1800 800
rect 1750 515 1765 785
rect 1785 515 1800 785
rect 1750 500 1800 515
rect 1850 785 1900 800
rect 1850 515 1865 785
rect 1885 515 1900 785
rect 1850 500 1900 515
rect 1950 785 2000 800
rect 1950 515 1965 785
rect 1985 515 2000 785
rect 1950 500 2000 515
rect 2050 785 2100 800
rect 2050 515 2065 785
rect 2085 515 2100 785
rect 2050 500 2100 515
rect 2150 785 2200 800
rect 2250 785 2300 800
rect 2150 515 2165 785
rect 2185 515 2200 785
rect 2250 515 2265 785
rect 2285 515 2300 785
rect 2150 500 2200 515
rect 2250 500 2300 515
rect 2350 785 2400 800
rect 2350 515 2365 785
rect 2385 515 2400 785
rect 2350 500 2400 515
rect 2450 785 2500 800
rect 2450 515 2465 785
rect 2485 515 2500 785
rect 2450 500 2500 515
rect 2550 785 2600 800
rect 2550 515 2565 785
rect 2585 515 2600 785
rect 2550 500 2600 515
rect 2650 785 2700 800
rect 2650 515 2665 785
rect 2685 515 2700 785
rect 2650 500 2700 515
rect 2750 785 2800 800
rect 2750 515 2765 785
rect 2785 515 2800 785
rect 2750 500 2800 515
rect 2850 785 2900 800
rect 2850 515 2865 785
rect 2885 515 2900 785
rect 2850 500 2900 515
rect -50 285 0 300
rect -50 15 -35 285
rect -15 15 0 285
rect -50 0 0 15
rect 50 285 100 300
rect 50 15 65 285
rect 85 15 100 285
rect 50 0 100 15
rect 150 285 200 300
rect 150 15 165 285
rect 185 15 200 285
rect 150 0 200 15
rect 250 285 300 300
rect 250 15 265 285
rect 285 15 300 285
rect 250 0 300 15
rect 350 285 400 300
rect 350 15 365 285
rect 385 15 400 285
rect 350 0 400 15
rect 450 285 500 300
rect 450 15 465 285
rect 485 15 500 285
rect 450 0 500 15
rect 550 285 600 300
rect 655 285 700 300
rect 550 15 565 285
rect 585 15 600 285
rect 655 15 670 285
rect 690 15 700 285
rect 550 0 600 15
rect 655 0 700 15
rect 750 285 800 300
rect 750 15 765 285
rect 785 15 800 285
rect 750 0 800 15
rect 850 0 875 300
rect 925 0 950 300
rect 1000 0 1025 300
rect 1075 0 1100 300
rect 1150 0 1175 300
rect 1225 0 1250 300
rect 1300 0 1325 300
rect 1375 0 1400 300
rect 1450 0 1475 300
rect 1525 0 1550 300
rect 1600 0 1625 300
rect 1675 0 1700 300
rect 1750 0 1775 300
rect 1825 0 1850 300
rect 1900 0 1925 300
rect 1975 0 2000 300
rect 2050 0 2075 300
rect 2125 0 2150 300
rect 2200 0 2225 300
rect 2275 285 2325 300
rect 2275 15 2290 285
rect 2310 15 2325 285
rect 2275 0 2325 15
rect 2375 285 2425 300
rect 2475 285 2525 300
rect 2375 15 2390 285
rect 2410 15 2425 285
rect 2475 15 2490 285
rect 2510 15 2525 285
rect 2375 0 2425 15
rect 2475 0 2525 15
rect 2575 285 2625 300
rect 2575 15 2590 285
rect 2610 15 2625 285
rect 2575 0 2625 15
rect 2675 285 2725 300
rect 2675 15 2690 285
rect 2710 15 2725 285
rect 2675 0 2725 15
rect 2775 285 2825 300
rect 2775 15 2790 285
rect 2810 15 2825 285
rect 2775 0 2825 15
rect 2875 285 2925 300
rect 2875 15 2890 285
rect 2910 15 2925 285
rect 2875 0 2925 15
rect 2975 285 3025 300
rect 2975 15 2990 285
rect 3010 15 3025 285
rect 2975 0 3025 15
rect 3075 285 3125 300
rect 3075 15 3090 285
rect 3110 15 3125 285
rect 3075 0 3125 15
<< pdiff >>
rect -50 1785 0 1800
rect -50 1515 -35 1785
rect -15 1515 0 1785
rect -50 1500 0 1515
rect 50 1785 100 1800
rect 50 1515 65 1785
rect 85 1515 100 1785
rect 50 1500 100 1515
rect 150 1785 200 1800
rect 150 1515 165 1785
rect 185 1515 200 1785
rect 150 1500 200 1515
rect 250 1785 300 1800
rect 250 1515 265 1785
rect 285 1515 300 1785
rect 250 1500 300 1515
rect 350 1785 400 1800
rect 350 1515 365 1785
rect 385 1515 400 1785
rect 350 1500 400 1515
rect 450 1785 500 1800
rect 450 1515 465 1785
rect 485 1515 500 1785
rect 450 1500 500 1515
rect 550 1785 600 1800
rect 655 1785 700 1800
rect 550 1515 565 1785
rect 585 1515 600 1785
rect 655 1515 670 1785
rect 690 1515 700 1785
rect 550 1500 600 1515
rect 655 1500 700 1515
rect 750 1785 800 1800
rect 750 1515 765 1785
rect 785 1515 800 1785
rect 750 1500 800 1515
rect 850 1500 875 1800
rect 925 1500 950 1800
rect 1000 1500 1025 1800
rect 1075 1500 1100 1800
rect 1150 1500 1175 1800
rect 1225 1500 1250 1800
rect 1300 1500 1325 1800
rect 1375 1500 1400 1800
rect 1450 1500 1475 1800
rect 1525 1500 1550 1800
rect 1600 1500 1625 1800
rect 1675 1500 1700 1800
rect 1750 1500 1775 1800
rect 1825 1500 1850 1800
rect 1900 1500 1925 1800
rect 1975 1500 2000 1800
rect 2050 1500 2075 1800
rect 2125 1500 2150 1800
rect 2200 1500 2225 1800
rect 2275 1785 2325 1800
rect 2275 1515 2290 1785
rect 2310 1515 2325 1785
rect 2275 1500 2325 1515
rect 2375 1785 2425 1800
rect 2475 1785 2525 1800
rect 2375 1515 2390 1785
rect 2410 1515 2425 1785
rect 2475 1515 2490 1785
rect 2510 1515 2525 1785
rect 2375 1500 2425 1515
rect 2475 1500 2525 1515
rect 2575 1785 2625 1800
rect 2575 1515 2590 1785
rect 2610 1515 2625 1785
rect 2575 1500 2625 1515
rect 2675 1785 2725 1800
rect 2675 1515 2690 1785
rect 2710 1515 2725 1785
rect 2675 1500 2725 1515
rect 2775 1785 2825 1800
rect 2775 1515 2790 1785
rect 2810 1515 2825 1785
rect 2775 1500 2825 1515
rect 2875 1785 2925 1800
rect 2875 1515 2890 1785
rect 2910 1515 2925 1785
rect 2875 1500 2925 1515
rect 2975 1785 3025 1800
rect 2975 1515 2990 1785
rect 3010 1515 3025 1785
rect 2975 1500 3025 1515
rect 3075 1785 3125 1800
rect 3075 1515 3090 1785
rect 3110 1515 3125 1785
rect 3075 1500 3125 1515
rect -250 1285 -200 1300
rect -250 1015 -235 1285
rect -215 1015 -200 1285
rect -250 1000 -200 1015
rect -150 1285 -100 1300
rect -150 1015 -135 1285
rect -115 1015 -100 1285
rect -150 1000 -100 1015
rect -50 1285 0 1300
rect -50 1015 -35 1285
rect -15 1015 0 1285
rect -50 1000 0 1015
rect 50 1285 100 1300
rect 50 1015 65 1285
rect 85 1015 100 1285
rect 50 1000 100 1015
rect 150 1285 200 1300
rect 150 1015 165 1285
rect 185 1015 200 1285
rect 150 1000 200 1015
rect 250 1285 300 1300
rect 250 1015 265 1285
rect 285 1015 300 1285
rect 250 1000 300 1015
rect 350 1285 400 1300
rect 455 1285 500 1300
rect 350 1015 365 1285
rect 390 1015 400 1285
rect 455 1015 470 1285
rect 490 1015 500 1285
rect 350 1000 400 1015
rect 455 1000 500 1015
rect 550 1285 600 1300
rect 550 1015 565 1285
rect 585 1015 600 1285
rect 550 1000 600 1015
rect 650 1285 700 1300
rect 650 1015 665 1285
rect 685 1015 700 1285
rect 650 1000 700 1015
rect 750 1285 800 1300
rect 750 1015 765 1285
rect 785 1015 800 1285
rect 750 1000 800 1015
rect 850 1285 900 1300
rect 850 1015 865 1285
rect 885 1015 900 1285
rect 850 1000 900 1015
rect 950 1285 1000 1300
rect 950 1015 965 1285
rect 985 1015 1000 1285
rect 950 1000 1000 1015
rect 1050 1285 1100 1300
rect 1050 1015 1065 1285
rect 1085 1015 1100 1285
rect 1050 1000 1100 1015
rect 1150 1285 1200 1300
rect 1150 1015 1165 1285
rect 1185 1015 1200 1285
rect 1150 1000 1200 1015
rect 1250 1285 1300 1300
rect 1250 1015 1265 1285
rect 1285 1015 1300 1285
rect 1250 1000 1300 1015
rect 1350 1285 1400 1300
rect 1350 1015 1365 1285
rect 1385 1015 1400 1285
rect 1350 1000 1400 1015
rect 1450 1285 1500 1300
rect 1450 1015 1465 1285
rect 1485 1015 1500 1285
rect 1450 1000 1500 1015
rect 1550 1285 1600 1300
rect 1550 1015 1565 1285
rect 1585 1015 1600 1285
rect 1550 1000 1600 1015
rect 1650 1285 1700 1300
rect 1650 1015 1665 1285
rect 1685 1015 1700 1285
rect 1650 1000 1700 1015
rect 1750 1285 1800 1300
rect 1750 1015 1765 1285
rect 1785 1015 1800 1285
rect 1750 1000 1800 1015
rect 1850 1285 1900 1300
rect 1850 1015 1865 1285
rect 1885 1015 1900 1285
rect 1850 1000 1900 1015
rect 1950 1285 2000 1300
rect 1950 1015 1965 1285
rect 1985 1015 2000 1285
rect 1950 1000 2000 1015
rect 2050 1285 2100 1300
rect 2050 1015 2065 1285
rect 2085 1015 2100 1285
rect 2050 1000 2100 1015
rect 2150 1285 2200 1300
rect 2150 1015 2165 1285
rect 2185 1015 2200 1285
rect 2150 1000 2200 1015
rect 2250 1285 2300 1300
rect 2250 1015 2265 1285
rect 2285 1015 2300 1285
rect 2250 1000 2300 1015
rect 2350 1285 2400 1300
rect 2350 1015 2365 1285
rect 2385 1015 2400 1285
rect 2350 1000 2400 1015
rect 2450 1285 2500 1300
rect 2450 1015 2465 1285
rect 2485 1015 2500 1285
rect 2450 1000 2500 1015
rect 2550 1285 2600 1300
rect 2550 1015 2565 1285
rect 2585 1015 2600 1285
rect 2550 1000 2600 1015
rect 2650 1295 2700 1300
rect 2650 1285 2695 1295
rect 2750 1285 2800 1300
rect 2650 1015 2665 1285
rect 2685 1015 2695 1285
rect 2750 1015 2765 1285
rect 2785 1015 2800 1285
rect 2650 1005 2695 1015
rect 2650 1000 2700 1005
rect 2750 1000 2800 1015
rect 2850 1285 2900 1300
rect 2850 1015 2865 1285
rect 2885 1015 2900 1285
rect 2850 1000 2900 1015
rect 2950 1285 3000 1300
rect 2950 1015 2965 1285
rect 2985 1015 3000 1285
rect 2950 1000 3000 1015
rect 3050 1285 3100 1300
rect 3050 1015 3065 1285
rect 3085 1015 3100 1285
rect 3050 1000 3100 1015
rect 3150 1285 3200 1300
rect 3150 1015 3165 1285
rect 3185 1015 3200 1285
rect 3150 1000 3200 1015
rect 3250 1285 3300 1300
rect 3250 1015 3265 1285
rect 3285 1015 3300 1285
rect 3250 1000 3300 1015
rect 3350 1295 3400 1300
rect 3350 1285 3390 1295
rect 3350 1015 3365 1285
rect 3385 1015 3390 1285
rect 3350 1005 3390 1015
rect 3350 1000 3400 1005
<< ndiffc >>
rect -35 515 -15 785
rect 65 515 85 785
rect 165 515 185 785
rect 265 515 285 785
rect 365 515 385 785
rect 465 515 485 785
rect 565 515 585 785
rect 665 515 685 785
rect 765 515 785 785
rect 865 515 885 785
rect 965 515 985 785
rect 1065 515 1085 785
rect 1165 515 1185 785
rect 1265 515 1285 785
rect 1365 515 1385 785
rect 1465 515 1485 785
rect 1565 515 1585 785
rect 1665 515 1685 785
rect 1765 515 1785 785
rect 1865 515 1885 785
rect 1965 515 1985 785
rect 2065 515 2085 785
rect 2165 515 2185 785
rect 2265 515 2285 785
rect 2365 515 2385 785
rect 2465 515 2485 785
rect 2565 515 2585 785
rect 2665 515 2685 785
rect 2765 515 2785 785
rect 2865 515 2885 785
rect -35 15 -15 285
rect 65 15 85 285
rect 165 15 185 285
rect 265 15 285 285
rect 365 15 385 285
rect 465 15 485 285
rect 565 15 585 285
rect 670 15 690 285
rect 765 15 785 285
rect 2290 15 2310 285
rect 2390 15 2410 285
rect 2490 15 2510 285
rect 2590 15 2610 285
rect 2690 15 2710 285
rect 2790 15 2810 285
rect 2890 15 2910 285
rect 2990 15 3010 285
rect 3090 15 3110 285
<< pdiffc >>
rect -35 1515 -15 1785
rect 65 1515 85 1785
rect 165 1515 185 1785
rect 265 1515 285 1785
rect 365 1515 385 1785
rect 465 1515 485 1785
rect 565 1515 585 1785
rect 670 1515 690 1785
rect 765 1515 785 1785
rect 2290 1515 2310 1785
rect 2390 1515 2410 1785
rect 2490 1515 2510 1785
rect 2590 1515 2610 1785
rect 2690 1515 2710 1785
rect 2790 1515 2810 1785
rect 2890 1515 2910 1785
rect 2990 1515 3010 1785
rect 3090 1515 3110 1785
rect -235 1015 -215 1285
rect -135 1015 -115 1285
rect -35 1015 -15 1285
rect 65 1015 85 1285
rect 165 1015 185 1285
rect 265 1015 285 1285
rect 365 1015 390 1285
rect 470 1015 490 1285
rect 565 1015 585 1285
rect 665 1015 685 1285
rect 765 1015 785 1285
rect 865 1015 885 1285
rect 965 1015 985 1285
rect 1065 1015 1085 1285
rect 1165 1015 1185 1285
rect 1265 1015 1285 1285
rect 1365 1015 1385 1285
rect 1465 1015 1485 1285
rect 1565 1015 1585 1285
rect 1665 1015 1685 1285
rect 1765 1015 1785 1285
rect 1865 1015 1885 1285
rect 1965 1015 1985 1285
rect 2065 1015 2085 1285
rect 2165 1015 2185 1285
rect 2265 1015 2285 1285
rect 2365 1015 2385 1285
rect 2465 1015 2485 1285
rect 2565 1015 2585 1285
rect 2665 1015 2685 1285
rect 2765 1015 2785 1285
rect 2865 1015 2885 1285
rect 2965 1015 2985 1285
rect 3065 1015 3085 1285
rect 3165 1015 3185 1285
rect 3265 1015 3285 1285
rect 3365 1015 3385 1285
<< psubdiff >>
rect -100 785 -50 800
rect -100 515 -85 785
rect -60 515 -50 785
rect -100 500 -50 515
rect 2200 785 2250 800
rect 2200 515 2215 785
rect 2235 515 2250 785
rect 2200 500 2250 515
rect 2900 785 2950 800
rect 2900 515 2915 785
rect 2935 515 2950 785
rect 2900 500 2950 515
rect -100 285 -50 300
rect -100 15 -85 285
rect -60 15 -50 285
rect -100 0 -50 15
rect 600 285 655 300
rect 600 15 615 285
rect 640 15 655 285
rect 600 0 655 15
rect 2425 285 2475 300
rect 2425 15 2440 285
rect 2460 15 2475 285
rect 2425 0 2475 15
rect 3125 285 3175 300
rect 3125 15 3140 285
rect 3160 15 3175 285
rect 3125 0 3175 15
<< nsubdiff >>
rect -100 1785 -50 1800
rect -100 1515 -85 1785
rect -65 1515 -50 1785
rect -100 1500 -50 1515
rect 600 1785 655 1800
rect 600 1515 615 1785
rect 640 1515 655 1785
rect 600 1500 655 1515
rect 2425 1785 2475 1800
rect 2425 1515 2440 1785
rect 2460 1515 2475 1785
rect 2425 1500 2475 1515
rect 3125 1785 3175 1800
rect 3125 1515 3140 1785
rect 3160 1515 3175 1785
rect 3125 1500 3175 1515
rect -300 1285 -250 1300
rect -300 1015 -285 1285
rect -260 1015 -250 1285
rect -300 1000 -250 1015
rect 400 1285 455 1300
rect 400 1015 415 1285
rect 440 1015 455 1285
rect 400 1000 455 1015
rect 2700 1295 2750 1300
rect 2695 1285 2750 1295
rect 2695 1015 2710 1285
rect 2735 1015 2750 1285
rect 2695 1005 2750 1015
rect 2700 1000 2750 1005
rect 3400 1295 3450 1300
rect 3390 1285 3450 1295
rect 3390 1015 3415 1285
rect 3435 1015 3450 1285
rect 3390 1005 3450 1015
rect 3400 1000 3450 1005
<< psubdiffcont >>
rect -85 515 -60 785
rect 2215 515 2235 785
rect 2915 515 2935 785
rect -85 15 -60 285
rect 615 15 640 285
rect 2440 15 2460 285
rect 3140 15 3160 285
<< nsubdiffcont >>
rect -85 1515 -65 1785
rect 615 1515 640 1785
rect 2440 1515 2460 1785
rect 3140 1515 3160 1785
rect -285 1015 -260 1285
rect 415 1015 440 1285
rect 2710 1015 2735 1285
rect 3415 1015 3435 1285
<< poly >>
rect 105 1855 145 1865
rect -45 1845 -5 1855
rect -45 1825 -35 1845
rect -15 1830 -5 1845
rect 100 1835 115 1855
rect 135 1840 2975 1855
rect 135 1835 150 1840
rect -15 1825 50 1830
rect -45 1815 50 1825
rect 0 1800 50 1815
rect 100 1800 150 1835
rect 200 1800 250 1840
rect 300 1800 350 1840
rect 400 1800 450 1840
rect 500 1800 550 1815
rect 700 1800 750 1815
rect 800 1800 850 1840
rect 875 1800 925 1840
rect 950 1800 1000 1840
rect 1025 1800 1075 1840
rect 1100 1800 1150 1840
rect 1175 1800 1225 1840
rect 1250 1800 1300 1840
rect 1325 1800 1375 1840
rect 1400 1800 1450 1840
rect 1475 1800 1525 1840
rect 1550 1800 1600 1840
rect 1625 1800 1675 1840
rect 1700 1800 1750 1840
rect 1775 1800 1825 1840
rect 1850 1800 1900 1840
rect 1925 1800 1975 1840
rect 2000 1800 2050 1840
rect 2075 1800 2125 1840
rect 2150 1800 2200 1840
rect 2225 1800 2275 1840
rect 2325 1800 2375 1815
rect 2525 1800 2575 1815
rect 2625 1800 2675 1840
rect 2725 1800 2775 1840
rect 2825 1800 2875 1840
rect 2925 1800 2975 1840
rect 3080 1845 3120 1855
rect 3080 1830 3090 1845
rect 3025 1825 3090 1830
rect 3110 1825 3120 1845
rect 3025 1815 3120 1825
rect 3025 1800 3075 1815
rect 0 1485 50 1500
rect 100 1405 150 1500
rect 200 1485 250 1500
rect 300 1485 350 1500
rect 400 1485 450 1500
rect 500 1485 550 1500
rect 700 1485 750 1500
rect 800 1485 850 1500
rect 875 1485 925 1500
rect 950 1485 1000 1500
rect 1025 1485 1075 1500
rect 1100 1485 1150 1500
rect 1175 1485 1225 1500
rect 1250 1485 1300 1500
rect 1325 1485 1375 1500
rect 1400 1485 1450 1500
rect 1475 1485 1525 1500
rect 1550 1485 1600 1500
rect 1625 1485 1675 1500
rect 1700 1485 1750 1500
rect 1775 1485 1825 1500
rect 1850 1485 1900 1500
rect 1925 1485 1975 1500
rect 2000 1485 2050 1500
rect 2075 1485 2125 1500
rect 2150 1485 2200 1500
rect 2225 1485 2275 1500
rect 2325 1485 2375 1500
rect 2525 1485 2575 1500
rect 2625 1485 2675 1500
rect 2725 1485 2775 1500
rect 2825 1485 2875 1500
rect 2925 1485 2975 1500
rect 3025 1485 3075 1500
rect 500 1475 750 1485
rect 500 1470 620 1475
rect 610 1455 620 1470
rect 640 1470 750 1475
rect 2325 1475 2575 1485
rect 2325 1470 2440 1475
rect 640 1455 650 1470
rect 610 1445 650 1455
rect 2430 1455 2440 1470
rect 2460 1470 2575 1475
rect 2460 1455 2470 1470
rect 2430 1445 2470 1455
rect 2880 1450 2920 1460
rect 2880 1430 2890 1450
rect 2910 1435 2920 1450
rect 2910 1430 3475 1435
rect 2880 1420 3475 1430
rect -320 1390 150 1405
rect -100 1385 100 1390
rect -245 1345 -205 1355
rect -245 1325 -235 1345
rect -215 1330 -205 1345
rect -100 1330 -50 1385
rect 3305 1345 3345 1355
rect -215 1325 -150 1330
rect -245 1315 -150 1325
rect -205 1310 -150 1315
rect -200 1300 -150 1310
rect -100 1315 250 1330
rect 600 1315 2550 1330
rect 3305 1325 3315 1345
rect 3335 1325 3345 1345
rect 3305 1315 3345 1325
rect -100 1300 -50 1315
rect 0 1300 50 1315
rect 100 1300 150 1315
rect 200 1300 250 1315
rect 300 1300 350 1315
rect 500 1300 550 1315
rect 600 1300 650 1315
rect 700 1300 750 1315
rect 800 1300 850 1315
rect 900 1300 950 1315
rect 1000 1300 1050 1315
rect 1100 1300 1150 1315
rect 1200 1300 1250 1315
rect 1300 1300 1350 1315
rect 1400 1300 1450 1315
rect 1500 1300 1550 1315
rect 1600 1300 1650 1315
rect 1700 1300 1750 1315
rect 1800 1300 1850 1315
rect 1900 1300 1950 1315
rect 2000 1300 2050 1315
rect 2100 1300 2150 1315
rect 2200 1300 2250 1315
rect 2300 1300 2350 1315
rect 2400 1300 2450 1315
rect 2500 1300 2550 1315
rect 2600 1300 2650 1315
rect 2800 1300 2850 1315
rect 2900 1300 2950 1315
rect 3000 1300 3050 1315
rect 3100 1300 3150 1315
rect 3200 1300 3250 1315
rect 3300 1300 3350 1315
rect -200 985 -150 1000
rect -100 985 -50 1000
rect 0 985 50 1000
rect 100 985 150 1000
rect 200 985 250 1000
rect 300 985 350 1000
rect 500 985 550 1000
rect 600 985 650 1000
rect 700 985 750 1000
rect 800 985 850 1000
rect 900 985 950 1000
rect 1000 985 1050 1000
rect 1100 985 1150 1000
rect 1200 985 1250 1000
rect 1300 985 1350 1000
rect 1400 985 1450 1000
rect 1500 985 1550 1000
rect 1600 985 1650 1000
rect 1700 985 1750 1000
rect 1800 985 1850 1000
rect 1900 985 1950 1000
rect 2000 985 2050 1000
rect 2100 985 2150 1000
rect 2200 985 2250 1000
rect 2300 985 2350 1000
rect 2400 985 2450 1000
rect 2500 985 2550 1000
rect 2600 985 2650 1000
rect 2800 985 2850 1000
rect 2900 985 2950 1000
rect 3000 985 3050 1000
rect 3100 985 3150 1000
rect 3200 985 3250 1000
rect 3300 985 3350 1000
rect 300 975 550 985
rect 300 970 420 975
rect -45 950 -5 960
rect -45 935 -35 950
rect -315 930 -35 935
rect -15 930 -5 950
rect 410 955 420 970
rect 440 970 550 975
rect 605 975 645 985
rect 440 955 450 970
rect 410 945 450 955
rect 605 955 615 975
rect 635 955 645 975
rect 2635 975 2815 985
rect 2635 970 2710 975
rect 605 945 645 955
rect 2700 955 2710 970
rect 2730 970 2815 975
rect 2900 975 3250 985
rect 2900 970 3215 975
rect 2730 955 2740 970
rect 2700 945 2740 955
rect 3205 955 3215 970
rect 3235 970 3250 975
rect 3235 955 3245 970
rect 3205 945 3245 955
rect -315 920 -5 930
rect -315 -40 -300 920
rect 605 895 620 945
rect 3460 895 3475 1420
rect -275 880 620 895
rect 2725 880 3475 895
rect -275 420 -260 880
rect 2725 860 2750 880
rect 105 845 145 855
rect 105 830 115 845
rect 100 825 115 830
rect 135 830 145 845
rect 2205 845 2245 855
rect 2205 830 2215 845
rect 135 825 2050 830
rect 100 815 2050 825
rect 2135 825 2215 830
rect 2235 830 2245 845
rect 2700 845 2750 860
rect 2700 830 2715 845
rect 2235 825 2315 830
rect 2135 815 2315 825
rect 2400 825 2715 830
rect 2735 825 2750 845
rect 2400 815 2750 825
rect 2805 845 2845 855
rect 2805 825 2815 845
rect 2835 825 2845 845
rect 2805 815 2845 825
rect 0 800 50 815
rect 100 800 150 815
rect 200 800 250 815
rect 300 800 350 815
rect 400 800 450 815
rect 500 800 550 815
rect 600 800 650 815
rect 700 800 750 815
rect 800 800 850 815
rect 900 800 950 815
rect 1000 800 1050 815
rect 1100 800 1150 815
rect 1200 800 1250 815
rect 1300 800 1350 815
rect 1400 800 1450 815
rect 1500 800 1550 815
rect 1600 800 1650 815
rect 1700 800 1750 815
rect 1800 800 1850 815
rect 1900 800 1950 815
rect 2000 800 2050 815
rect 2100 800 2150 815
rect 2300 800 2350 815
rect 2400 800 2450 815
rect 2500 800 2550 815
rect 2600 800 2650 815
rect 2700 800 2750 815
rect 2800 800 2850 815
rect 0 485 50 500
rect 100 485 150 500
rect 200 485 250 500
rect 300 485 350 500
rect 400 485 450 500
rect 500 485 550 500
rect 600 485 650 500
rect 700 485 750 500
rect 800 485 850 500
rect 900 485 950 500
rect 1000 485 1050 500
rect 1100 485 1150 500
rect 1200 485 1250 500
rect 1300 485 1350 500
rect 1400 485 1450 500
rect 1500 485 1550 500
rect 1600 485 1650 500
rect 1700 485 1750 500
rect 1800 485 1850 500
rect 1900 485 1950 500
rect 2000 485 2050 500
rect 2100 485 2150 500
rect 2300 485 2350 500
rect 2400 485 2450 500
rect 2500 485 2550 500
rect 2600 485 2650 500
rect 2700 485 2750 500
rect 2800 485 2850 500
rect -45 475 15 485
rect -45 455 -35 475
rect -15 470 15 475
rect -15 455 -5 470
rect -45 445 -5 455
rect -275 405 770 420
rect 755 380 770 405
rect 755 370 795 380
rect -45 345 -5 355
rect -45 325 -35 345
rect -15 330 -5 345
rect 610 345 650 355
rect 610 330 620 345
rect -15 325 20 330
rect -45 315 20 325
rect 535 325 620 330
rect 640 330 650 345
rect 755 350 765 370
rect 785 350 795 370
rect 755 340 795 350
rect 2430 345 2470 355
rect 2430 330 2440 345
rect 640 325 725 330
rect 535 315 725 325
rect 2360 325 2440 330
rect 2460 330 2470 345
rect 2460 325 2540 330
rect 2360 315 2540 325
rect 0 300 50 315
rect 100 300 150 315
rect 200 300 250 315
rect 300 300 350 315
rect 400 300 450 315
rect 500 300 550 315
rect 700 300 750 315
rect 800 300 850 315
rect 875 300 925 315
rect 950 300 1000 315
rect 1025 300 1075 315
rect 1100 300 1150 315
rect 1175 300 1225 315
rect 1250 300 1300 315
rect 1325 300 1375 315
rect 1400 300 1450 315
rect 1475 300 1525 315
rect 1550 300 1600 315
rect 1625 300 1675 315
rect 1700 300 1750 315
rect 1775 300 1825 315
rect 1850 300 1900 315
rect 1925 300 1975 315
rect 2000 300 2050 315
rect 2075 300 2125 315
rect 2150 300 2200 315
rect 2225 300 2275 315
rect 2325 300 2375 315
rect 2525 300 2575 315
rect 2625 300 2675 315
rect 2725 300 2775 315
rect 2825 300 2875 315
rect 2925 300 2975 315
rect 3025 300 3075 315
rect 0 -15 50 0
rect 100 -25 150 0
rect 100 -40 115 -25
rect -315 -45 115 -40
rect 135 -40 150 -25
rect 200 -40 250 0
rect 300 -40 350 0
rect 400 -40 450 0
rect 500 -15 550 0
rect 700 -15 750 0
rect 800 -40 850 0
rect 875 -40 925 0
rect 950 -40 1000 0
rect 1025 -40 1075 0
rect 1100 -40 1150 0
rect 1175 -40 1225 0
rect 1250 -40 1300 0
rect 1325 -40 1375 0
rect 1400 -40 1450 0
rect 1475 -40 1525 0
rect 1550 -40 1600 0
rect 1625 -40 1675 0
rect 1700 -40 1750 0
rect 1775 -40 1825 0
rect 1850 -40 1900 0
rect 1925 -40 1975 0
rect 2000 -40 2050 0
rect 2075 -40 2125 0
rect 2150 -40 2200 0
rect 2225 -40 2275 0
rect 2325 -15 2375 0
rect 2525 -15 2575 0
rect 2625 -40 2675 0
rect 2725 -40 2775 0
rect 2825 -40 2875 0
rect 2925 -40 2975 0
rect 3025 -15 3075 0
rect 3060 -25 3120 -15
rect 3060 -30 3090 -25
rect 135 -45 2975 -40
rect -315 -55 2975 -45
rect 3080 -45 3090 -30
rect 3110 -45 3120 -25
rect 3080 -55 3120 -45
<< polycont >>
rect -35 1825 -15 1845
rect 115 1835 135 1855
rect 3090 1825 3110 1845
rect 620 1455 640 1475
rect 2440 1455 2460 1475
rect 2890 1430 2910 1450
rect -235 1325 -215 1345
rect 3315 1325 3335 1345
rect -35 930 -15 950
rect 420 955 440 975
rect 615 955 635 975
rect 2710 955 2730 975
rect 3215 955 3235 975
rect 115 825 135 845
rect 2215 825 2235 845
rect 2715 825 2735 845
rect 2815 825 2835 845
rect -35 455 -15 475
rect -35 325 -15 345
rect 620 325 640 345
rect 765 350 785 370
rect 2440 325 2460 345
rect 115 -45 135 -25
rect 3090 -45 3110 -25
<< locali >>
rect 105 1855 145 1865
rect -45 1845 -5 1855
rect 105 1845 115 1855
rect -45 1825 -35 1845
rect -15 1825 -5 1845
rect -45 1795 -5 1825
rect -95 1785 -5 1795
rect -95 1515 -85 1785
rect -65 1515 -35 1785
rect -15 1515 -5 1785
rect -95 1505 -5 1515
rect 55 1835 115 1845
rect 135 1845 145 1855
rect 3080 1845 3120 1855
rect 135 1835 290 1845
rect 55 1825 290 1835
rect 55 1785 95 1825
rect 260 1795 290 1825
rect 3080 1825 3090 1845
rect 3110 1825 3120 1845
rect 3080 1795 3120 1825
rect 55 1515 65 1785
rect 85 1515 95 1785
rect 55 1505 95 1515
rect 155 1785 195 1795
rect 155 1515 165 1785
rect 185 1515 195 1785
rect 155 1505 195 1515
rect 255 1785 295 1795
rect 255 1515 265 1785
rect 285 1515 295 1785
rect 255 1505 295 1515
rect 355 1785 395 1795
rect 355 1515 365 1785
rect 385 1515 395 1785
rect 355 1505 395 1515
rect 455 1785 495 1795
rect 455 1515 465 1785
rect 485 1515 495 1785
rect 455 1505 495 1515
rect 555 1785 700 1795
rect 555 1515 565 1785
rect 585 1515 615 1785
rect 640 1515 670 1785
rect 690 1515 700 1785
rect 555 1505 700 1515
rect 755 1785 800 1795
rect 755 1515 765 1785
rect 785 1515 800 1785
rect 755 1505 800 1515
rect 2280 1785 2320 1795
rect 2280 1515 2290 1785
rect 2310 1515 2320 1785
rect 2280 1505 2320 1515
rect 2380 1785 2520 1795
rect 2380 1515 2390 1785
rect 2410 1515 2440 1785
rect 2460 1515 2490 1785
rect 2510 1515 2520 1785
rect 2380 1505 2520 1515
rect 2580 1785 2620 1795
rect 2580 1515 2590 1785
rect 2610 1515 2620 1785
rect 2580 1505 2620 1515
rect 2680 1785 2720 1795
rect 2680 1515 2690 1785
rect 2710 1515 2720 1785
rect 610 1475 650 1505
rect 610 1455 620 1475
rect 640 1455 650 1475
rect 610 1445 650 1455
rect 755 1395 775 1505
rect 2430 1475 2470 1505
rect 2430 1455 2440 1475
rect 2460 1455 2470 1475
rect 2680 1485 2720 1515
rect 2780 1785 2820 1795
rect 2780 1515 2790 1785
rect 2810 1515 2820 1785
rect 2780 1505 2820 1515
rect 2880 1785 2920 1795
rect 2880 1515 2890 1785
rect 2910 1515 2920 1785
rect 2880 1485 2920 1515
rect 2980 1785 3020 1795
rect 2980 1515 2990 1785
rect 3010 1515 3020 1785
rect 2980 1505 3020 1515
rect 3080 1785 3170 1795
rect 3080 1515 3090 1785
rect 3110 1515 3140 1785
rect 3160 1515 3170 1785
rect 3080 1505 3170 1515
rect 2680 1460 2920 1485
rect 2430 1445 2470 1455
rect 2880 1450 2920 1460
rect 2880 1430 2890 1450
rect 2910 1430 2920 1450
rect 2880 1420 2920 1430
rect -340 1375 775 1395
rect -340 855 -320 1375
rect -245 1345 -205 1355
rect -245 1325 -235 1345
rect -215 1325 -205 1345
rect 3305 1345 3345 1355
rect -245 1295 -205 1325
rect 655 1315 3195 1335
rect 3305 1325 3315 1345
rect 3335 1335 3345 1345
rect 3335 1325 3375 1335
rect 3305 1315 3375 1325
rect -295 1285 -205 1295
rect -295 1015 -285 1285
rect -260 1015 -235 1285
rect -215 1015 -205 1285
rect -295 1005 -205 1015
rect -145 1285 -105 1295
rect -145 1015 -135 1285
rect -115 1015 -105 1285
rect -145 1005 -105 1015
rect -45 1285 -5 1295
rect -45 1015 -35 1285
rect -15 1015 -5 1285
rect -45 985 -5 1015
rect 55 1285 95 1295
rect 55 1015 65 1285
rect 85 1015 95 1285
rect 55 1005 95 1015
rect 155 1285 195 1295
rect 155 1015 165 1285
rect 185 1015 195 1285
rect 155 985 195 1015
rect 255 1285 295 1295
rect 255 1015 265 1285
rect 285 1015 295 1285
rect 255 1005 295 1015
rect 355 1285 500 1295
rect 355 1015 365 1285
rect 390 1015 415 1285
rect 440 1015 470 1285
rect 490 1015 500 1285
rect 355 1005 500 1015
rect 555 1285 595 1295
rect 555 1015 565 1285
rect 585 1015 595 1285
rect 555 1005 595 1015
rect 655 1285 695 1315
rect 655 1015 665 1285
rect 685 1015 695 1285
rect 655 1005 695 1015
rect 755 1285 795 1295
rect 755 1015 765 1285
rect 785 1015 795 1285
rect -45 965 195 985
rect 410 975 450 1005
rect 755 985 795 1015
rect 855 1285 895 1315
rect 855 1015 865 1285
rect 885 1015 895 1285
rect 855 1005 895 1015
rect 955 1285 995 1295
rect 955 1015 965 1285
rect 985 1015 995 1285
rect 955 985 995 1015
rect 1055 1285 1095 1315
rect 1055 1015 1065 1285
rect 1085 1015 1095 1285
rect 1055 1005 1095 1015
rect 1155 1285 1195 1295
rect 1155 1015 1165 1285
rect 1185 1015 1195 1285
rect 1155 985 1195 1015
rect 1255 1285 1295 1315
rect 1255 1015 1265 1285
rect 1285 1015 1295 1285
rect 1255 1005 1295 1015
rect 1355 1285 1395 1295
rect 1355 1015 1365 1285
rect 1385 1015 1395 1285
rect 1355 985 1395 1015
rect 1455 1285 1495 1315
rect 1455 1015 1465 1285
rect 1485 1015 1495 1285
rect 1455 1005 1495 1015
rect 1555 1285 1595 1295
rect 1555 1015 1565 1285
rect 1585 1015 1595 1285
rect 1555 1005 1595 1015
rect 1655 1285 1695 1315
rect 1655 1015 1665 1285
rect 1685 1015 1695 1285
rect 1655 1005 1695 1015
rect 1755 1285 1795 1295
rect 1755 1015 1765 1285
rect 1785 1015 1795 1285
rect 1755 985 1795 1015
rect 1855 1285 1895 1315
rect 1855 1015 1865 1285
rect 1885 1015 1895 1285
rect 1855 1005 1895 1015
rect 1955 1285 1995 1295
rect 1955 1015 1965 1285
rect 1985 1015 1995 1285
rect 1955 985 1995 1015
rect 2055 1285 2095 1315
rect 2055 1015 2065 1285
rect 2085 1015 2095 1285
rect 2055 1005 2095 1015
rect 2155 1285 2195 1295
rect 2155 1015 2165 1285
rect 2185 1015 2195 1285
rect 2155 985 2195 1015
rect 2255 1285 2295 1315
rect 2255 1015 2265 1285
rect 2285 1015 2295 1285
rect 2255 1005 2295 1015
rect 2355 1285 2395 1295
rect 2355 1015 2365 1285
rect 2385 1015 2395 1285
rect 2355 985 2395 1015
rect 2455 1285 2495 1315
rect 2455 1015 2465 1285
rect 2485 1015 2495 1285
rect 2455 1005 2495 1015
rect 2555 1285 2595 1295
rect 2555 1015 2565 1285
rect 2585 1015 2595 1285
rect 2555 1005 2595 1015
rect 2655 1285 2795 1295
rect 2655 1015 2665 1285
rect 2685 1015 2710 1285
rect 2735 1015 2765 1285
rect 2785 1015 2795 1285
rect 2655 1005 2795 1015
rect 2855 1285 2895 1295
rect 2855 1015 2865 1285
rect 2885 1015 2895 1285
rect -45 950 -5 965
rect -45 930 -35 950
rect -15 930 -5 950
rect 410 955 420 975
rect 440 955 450 975
rect 410 945 450 955
rect 605 975 2395 985
rect 605 955 615 975
rect 635 965 2395 975
rect 2700 975 2740 1005
rect 635 955 645 965
rect 605 945 645 955
rect 2700 955 2710 975
rect 2730 955 2740 975
rect 2855 985 2895 1015
rect 2955 1285 2995 1315
rect 2955 1015 2965 1285
rect 2985 1015 2995 1285
rect 2955 1005 2995 1015
rect 3055 1285 3095 1295
rect 3055 1015 3065 1285
rect 3085 1015 3095 1285
rect 3055 985 3095 1015
rect 3155 1285 3195 1315
rect 3355 1295 3375 1315
rect 3155 1015 3165 1285
rect 3185 1015 3195 1285
rect 3155 1005 3195 1015
rect 3255 1285 3295 1295
rect 3255 1015 3265 1285
rect 3285 1015 3295 1285
rect 3255 985 3295 1015
rect 3355 1285 3445 1295
rect 3355 1015 3365 1285
rect 3385 1015 3415 1285
rect 3435 1015 3445 1285
rect 3355 1005 3445 1015
rect 2855 975 3295 985
rect 2855 965 3215 975
rect 2700 945 2740 955
rect -45 920 -5 930
rect -340 845 145 855
rect -340 835 115 845
rect 105 825 115 835
rect 135 835 145 845
rect 2205 845 2245 855
rect 135 825 1895 835
rect 105 815 1895 825
rect -95 785 -5 795
rect -95 515 -85 785
rect -60 515 -35 785
rect -15 515 -5 785
rect -95 505 -5 515
rect 55 785 95 795
rect 55 515 65 785
rect 85 515 95 785
rect 55 505 95 515
rect 155 785 195 795
rect 155 515 165 785
rect 185 515 195 785
rect -45 475 -5 505
rect -45 455 -35 475
rect -15 455 -5 475
rect 155 485 195 515
rect 255 785 295 815
rect 255 515 265 785
rect 285 515 295 785
rect 255 505 295 515
rect 355 785 395 795
rect 355 515 365 785
rect 385 515 395 785
rect 355 485 395 515
rect 455 785 495 815
rect 455 515 465 785
rect 485 515 495 785
rect 455 505 495 515
rect 555 785 595 795
rect 555 515 565 785
rect 585 515 595 785
rect 555 485 595 515
rect 655 785 695 815
rect 655 515 665 785
rect 685 515 695 785
rect 655 505 695 515
rect 755 785 795 795
rect 755 515 765 785
rect 785 515 795 785
rect 755 485 795 515
rect 855 785 895 815
rect 855 515 865 785
rect 885 515 895 785
rect 855 505 895 515
rect 955 785 995 795
rect 955 515 965 785
rect 985 515 995 785
rect 955 485 995 515
rect 1055 785 1095 795
rect 1055 515 1065 785
rect 1085 515 1095 785
rect 1055 505 1095 515
rect 1155 785 1195 795
rect 1155 515 1165 785
rect 1185 515 1195 785
rect 1155 485 1195 515
rect 1255 785 1295 815
rect 1255 515 1265 785
rect 1285 515 1295 785
rect 1255 505 1295 515
rect 1355 785 1395 795
rect 1355 515 1365 785
rect 1385 515 1395 785
rect 1355 485 1395 515
rect 1455 785 1495 815
rect 1455 515 1465 785
rect 1485 515 1495 785
rect 1455 505 1495 515
rect 1555 785 1595 795
rect 1555 515 1565 785
rect 1585 515 1595 785
rect 1555 485 1595 515
rect 1655 785 1695 815
rect 1655 515 1665 785
rect 1685 515 1695 785
rect 1655 505 1695 515
rect 1755 785 1795 795
rect 1755 515 1765 785
rect 1785 515 1795 785
rect 1755 485 1795 515
rect 1855 785 1895 815
rect 2205 825 2215 845
rect 2235 825 2245 845
rect 2705 845 2745 855
rect 2705 835 2715 845
rect 2205 795 2245 825
rect 2455 825 2715 835
rect 2735 825 2745 845
rect 2455 815 2745 825
rect 2805 845 2845 855
rect 2805 825 2815 845
rect 2835 835 2845 845
rect 2835 825 2875 835
rect 2805 815 2875 825
rect 1855 515 1865 785
rect 1885 515 1895 785
rect 1855 505 1895 515
rect 1955 785 1995 795
rect 1955 515 1965 785
rect 1985 515 1995 785
rect 1955 485 1995 515
rect 2055 785 2095 795
rect 2055 515 2065 785
rect 2085 515 2095 785
rect 2055 505 2095 515
rect 2155 785 2295 795
rect 2155 515 2165 785
rect 2185 515 2215 785
rect 2235 515 2265 785
rect 2285 515 2295 785
rect 2155 505 2295 515
rect 2355 785 2395 795
rect 2355 515 2365 785
rect 2385 515 2395 785
rect 2355 485 2395 515
rect 2455 785 2495 815
rect 2455 515 2465 785
rect 2485 515 2495 785
rect 2455 505 2495 515
rect 2555 785 2595 795
rect 2555 515 2565 785
rect 2585 515 2595 785
rect 2555 485 2595 515
rect 2655 785 2695 815
rect 2855 795 2875 815
rect 2655 515 2665 785
rect 2685 515 2695 785
rect 2655 505 2695 515
rect 2755 785 2795 795
rect 2755 515 2765 785
rect 2785 515 2795 785
rect 2755 485 2795 515
rect 2855 785 2945 795
rect 2855 515 2865 785
rect 2885 515 2915 785
rect 2935 515 2945 785
rect 2855 505 2945 515
rect 155 465 2795 485
rect -45 445 -5 455
rect 755 370 795 380
rect -45 345 -5 355
rect -45 325 -35 345
rect -15 325 -5 345
rect -45 295 -5 325
rect 610 345 650 355
rect 610 325 620 345
rect 640 325 650 345
rect 610 295 650 325
rect 755 350 765 370
rect 785 350 795 370
rect 3055 355 3075 965
rect 3205 955 3215 965
rect 3235 965 3295 975
rect 3235 955 3475 965
rect 3205 945 3475 955
rect 755 295 795 350
rect 2430 345 2470 355
rect 2430 325 2440 345
rect 2460 325 2470 345
rect 2900 335 3075 355
rect 2430 295 2470 325
rect 2680 315 2920 335
rect -95 285 -5 295
rect -95 15 -85 285
rect -60 15 -35 285
rect -15 15 -5 285
rect -95 5 -5 15
rect 55 285 95 295
rect 55 15 65 285
rect 85 15 95 285
rect 55 5 95 15
rect 155 285 195 295
rect 155 15 165 285
rect 185 15 195 285
rect 155 -15 195 15
rect 255 285 295 295
rect 255 15 265 285
rect 285 15 295 285
rect 255 5 295 15
rect 355 285 395 295
rect 355 15 365 285
rect 385 15 395 285
rect 355 -15 395 15
rect 455 285 495 295
rect 455 15 465 285
rect 485 15 495 285
rect 455 5 495 15
rect 555 285 700 295
rect 555 15 565 285
rect 585 15 615 285
rect 640 15 670 285
rect 690 15 700 285
rect 555 5 700 15
rect 755 285 800 295
rect 755 15 765 285
rect 785 15 800 285
rect 755 5 800 15
rect 2280 285 2320 295
rect 2280 15 2290 285
rect 2310 15 2320 285
rect 2280 5 2320 15
rect 2380 285 2520 295
rect 2380 15 2390 285
rect 2410 15 2440 285
rect 2460 15 2490 285
rect 2510 15 2520 285
rect 2380 5 2520 15
rect 2580 285 2620 295
rect 2580 15 2590 285
rect 2610 15 2620 285
rect 2580 5 2620 15
rect 2680 285 2720 315
rect 2680 15 2690 285
rect 2710 15 2720 285
rect 2680 5 2720 15
rect 2780 285 2820 295
rect 2780 15 2790 285
rect 2810 15 2820 285
rect 2780 5 2820 15
rect 2880 285 2920 315
rect 2880 15 2890 285
rect 2910 15 2920 285
rect 2880 5 2920 15
rect 2980 285 3020 295
rect 2980 15 2990 285
rect 3010 15 3020 285
rect 2980 5 3020 15
rect 3080 285 3170 295
rect 3080 15 3090 285
rect 3110 15 3140 285
rect 3160 15 3170 285
rect 3080 5 3170 15
rect 105 -25 395 -15
rect 105 -45 115 -25
rect 135 -35 395 -25
rect 3080 -25 3120 5
rect 135 -45 145 -35
rect 105 -55 145 -45
rect 3080 -45 3090 -25
rect 3110 -45 3120 -25
rect 3080 -55 3120 -45
<< viali >>
rect -85 1515 -65 1785
rect -35 1515 -15 1785
rect 165 1515 185 1785
rect 365 1515 385 1785
rect 565 1515 585 1785
rect 615 1515 640 1785
rect 670 1515 690 1785
rect 2290 1515 2310 1785
rect 2390 1515 2410 1785
rect 2440 1515 2460 1785
rect 2490 1515 2510 1785
rect 2590 1515 2610 1785
rect 2790 1515 2810 1785
rect 2990 1515 3010 1785
rect 3090 1515 3110 1785
rect 3140 1515 3160 1785
rect -285 1015 -260 1285
rect -235 1015 -215 1285
rect -135 1015 -115 1285
rect 65 1015 85 1285
rect 265 1015 285 1285
rect 365 1015 390 1285
rect 415 1015 440 1285
rect 470 1015 490 1285
rect 565 1015 585 1285
rect 1565 1015 1585 1285
rect 2565 1015 2585 1285
rect 2665 1015 2685 1285
rect 2710 1015 2735 1285
rect 2765 1015 2785 1285
rect 3365 1015 3385 1285
rect 3415 1015 3435 1285
rect -85 515 -60 785
rect -35 515 -15 785
rect 65 515 85 785
rect 1065 515 1085 785
rect 2065 515 2085 785
rect 2165 515 2185 785
rect 2215 515 2235 785
rect 2265 515 2285 785
rect 2865 515 2885 785
rect 2915 515 2935 785
rect -85 15 -60 285
rect -35 15 -15 285
rect 65 15 85 285
rect 265 15 285 285
rect 465 15 485 285
rect 565 15 585 285
rect 615 15 640 285
rect 670 15 690 285
rect 2290 15 2310 285
rect 2390 15 2410 285
rect 2440 15 2460 285
rect 2490 15 2510 285
rect 2590 15 2610 285
rect 2790 15 2810 285
rect 2990 15 3010 285
rect 3090 15 3110 285
rect 3140 15 3160 285
<< metal1 >>
rect -320 1785 3455 1800
rect -320 1515 -85 1785
rect -65 1515 -35 1785
rect -15 1515 165 1785
rect 185 1515 365 1785
rect 385 1515 565 1785
rect 585 1515 615 1785
rect 640 1515 670 1785
rect 690 1515 2290 1785
rect 2310 1515 2390 1785
rect 2410 1515 2440 1785
rect 2460 1515 2490 1785
rect 2510 1515 2590 1785
rect 2610 1515 2790 1785
rect 2810 1515 2990 1785
rect 3010 1515 3090 1785
rect 3110 1515 3140 1785
rect 3160 1515 3455 1785
rect -320 1285 3455 1515
rect -320 1015 -285 1285
rect -260 1015 -235 1285
rect -215 1015 -135 1285
rect -115 1015 65 1285
rect 85 1015 265 1285
rect 285 1015 365 1285
rect 390 1015 415 1285
rect 440 1015 470 1285
rect 490 1015 565 1285
rect 585 1015 1565 1285
rect 1585 1015 2565 1285
rect 2585 1015 2665 1285
rect 2685 1015 2710 1285
rect 2735 1015 2765 1285
rect 2785 1015 3365 1285
rect 3385 1015 3415 1285
rect 3435 1015 3455 1285
rect -320 1000 3455 1015
rect -120 785 3195 805
rect -120 515 -85 785
rect -60 515 -35 785
rect -15 515 65 785
rect 85 515 1065 785
rect 1085 515 2065 785
rect 2085 515 2165 785
rect 2185 515 2215 785
rect 2235 515 2265 785
rect 2285 515 2865 785
rect 2885 515 2915 785
rect 2935 515 3195 785
rect -120 285 3195 515
rect -120 15 -85 285
rect -60 15 -35 285
rect -15 15 65 285
rect 85 15 265 285
rect 285 15 465 285
rect 485 15 565 285
rect 585 15 615 285
rect 640 15 670 285
rect 690 15 2290 285
rect 2310 15 2390 285
rect 2410 15 2440 285
rect 2460 15 2490 285
rect 2510 15 2590 285
rect 2610 15 2790 285
rect 2810 15 2990 285
rect 3010 15 3090 285
rect 3110 15 3140 285
rect 3160 15 3195 285
rect -120 0 3195 15
<< labels >>
rlabel metal1 -320 1420 -320 1420 7 VP
port 1 w
rlabel metal1 -120 305 -120 305 7 VN
port 2 w
rlabel poly -320 1395 -320 1395 7 Vbp
port 3 w
rlabel poly -315 -50 -315 -50 7 Vbn
port 4 w
rlabel locali 3475 955 3475 955 3 Vcp
port 6 e
rlabel locali 680 1305 680 1305 7 net42
rlabel pdiff 860 1700 860 1700 7 net1
rlabel locali 870 810 870 810 7 net39
rlabel locali 165 485 165 485 7 net40
rlabel pdiff 2210 1580 2210 1580 7 net19
<< end >>
