magic
tech sky130A
timestamp 1614784726
<< nwell >>
rect -85 415 435 745
<< nmos >>
rect 0 225 15 325
rect 40 225 55 325
rect 235 245 250 345
rect 300 245 315 345
rect -20 -10 -5 90
rect 20 -10 35 90
rect 235 -10 250 90
rect 300 -10 315 90
<< pmos >>
rect 0 625 15 725
rect 40 625 55 725
rect 235 625 250 725
rect 275 625 290 725
rect 0 435 15 535
rect 65 435 80 535
rect 235 435 250 535
rect 275 435 290 535
<< ndiff >>
rect -50 310 0 325
rect -50 240 -35 310
rect -15 240 0 310
rect -50 225 0 240
rect 15 225 40 325
rect 55 310 105 325
rect 55 240 70 310
rect 90 240 105 310
rect 55 225 105 240
rect 185 330 235 345
rect 185 260 200 330
rect 220 260 235 330
rect 185 245 235 260
rect 250 330 300 345
rect 250 260 265 330
rect 285 260 300 330
rect 250 245 300 260
rect 315 330 365 345
rect 315 260 330 330
rect 350 260 365 330
rect 315 245 365 260
rect -70 75 -20 90
rect -70 5 -55 75
rect -35 5 -20 75
rect -70 -10 -20 5
rect -5 -10 20 90
rect 35 75 85 90
rect 35 5 50 75
rect 70 5 85 75
rect 35 -10 85 5
rect 185 75 235 90
rect 185 5 200 75
rect 220 5 235 75
rect 185 -10 235 5
rect 250 75 300 90
rect 250 5 265 75
rect 285 5 300 75
rect 250 -10 300 5
rect 315 75 365 90
rect 315 5 330 75
rect 350 5 365 75
rect 315 -10 365 5
<< pdiff >>
rect -50 710 0 725
rect -50 640 -35 710
rect -15 640 0 710
rect -50 625 0 640
rect 15 625 40 725
rect 55 710 105 725
rect 55 640 70 710
rect 90 640 105 710
rect 55 625 105 640
rect 185 710 235 725
rect 185 640 200 710
rect 220 640 235 710
rect 185 625 235 640
rect 250 625 275 725
rect 290 710 340 725
rect 290 640 305 710
rect 325 640 340 710
rect 290 625 340 640
rect -50 520 0 535
rect -50 450 -35 520
rect -15 450 0 520
rect -50 435 0 450
rect 15 520 65 535
rect 15 450 30 520
rect 50 450 65 520
rect 15 435 65 450
rect 80 520 130 535
rect 80 450 95 520
rect 115 450 130 520
rect 80 435 130 450
rect 185 520 235 535
rect 185 450 200 520
rect 220 450 235 520
rect 185 435 235 450
rect 250 435 275 535
rect 290 520 340 535
rect 290 450 305 520
rect 325 450 340 520
rect 290 435 340 450
<< ndiffc >>
rect -35 240 -15 310
rect 70 240 90 310
rect 200 260 220 330
rect 265 260 285 330
rect 330 260 350 330
rect -55 5 -35 75
rect 50 5 70 75
rect 200 5 220 75
rect 265 5 285 75
rect 330 5 350 75
<< pdiffc >>
rect -35 640 -15 710
rect 70 640 90 710
rect 200 640 220 710
rect 305 640 325 710
rect -35 450 -15 520
rect 30 450 50 520
rect 95 450 115 520
rect 200 450 220 520
rect 305 450 325 520
<< psubdiff >>
rect 85 75 135 90
rect 85 5 100 75
rect 120 5 135 75
rect 85 -10 135 5
rect 365 75 415 90
rect 365 5 380 75
rect 400 5 415 75
rect 365 -10 415 5
<< nsubdiff >>
rect 105 710 155 725
rect 105 640 120 710
rect 140 640 155 710
rect 105 625 155 640
rect 340 710 390 725
rect 340 640 355 710
rect 375 640 390 710
rect 340 625 390 640
<< psubdiffcont >>
rect 100 5 120 75
rect 380 5 400 75
<< nsubdiffcont >>
rect 120 640 140 710
rect 355 640 375 710
<< poly >>
rect 0 725 15 740
rect 40 725 55 740
rect 235 725 250 740
rect 275 725 290 740
rect 0 535 15 625
rect 40 600 55 625
rect 40 590 80 600
rect 40 570 50 590
rect 70 570 80 590
rect 40 560 80 570
rect 65 535 80 560
rect 235 535 250 625
rect 275 610 290 625
rect 275 595 380 610
rect 275 535 290 550
rect -65 405 -25 415
rect -65 400 -55 405
rect -85 385 -55 400
rect -35 385 -25 405
rect -65 375 -25 385
rect 0 325 15 435
rect 65 420 80 435
rect 65 405 135 420
rect 50 370 90 380
rect 50 355 60 370
rect 40 350 60 355
rect 80 350 90 370
rect 40 340 90 350
rect 40 325 55 340
rect 0 210 15 225
rect -20 195 15 210
rect -20 90 -5 195
rect 40 185 55 225
rect 120 185 135 405
rect 235 345 250 435
rect 275 420 290 435
rect 275 405 315 420
rect 300 345 315 405
rect 365 400 380 595
rect 340 390 435 400
rect 340 370 350 390
rect 370 385 435 390
rect 370 370 380 385
rect 340 360 380 370
rect 170 200 210 210
rect 170 185 180 200
rect 40 180 180 185
rect 200 180 210 200
rect 40 175 210 180
rect 40 160 65 175
rect 20 155 65 160
rect 85 170 210 175
rect 85 155 95 170
rect 20 145 95 155
rect 20 90 35 145
rect 235 90 250 245
rect 300 190 315 245
rect 340 220 380 230
rect 340 200 350 220
rect 370 200 380 220
rect 340 190 380 200
rect 275 180 315 190
rect 275 160 285 180
rect 305 160 315 180
rect 275 150 315 160
rect 365 120 380 190
rect 300 105 380 120
rect 300 90 315 105
rect -20 -40 -5 -10
rect 20 -25 35 -10
rect -45 -50 -5 -40
rect -45 -70 -35 -50
rect -15 -70 -5 -50
rect -45 -80 -5 -70
rect 235 -40 250 -10
rect 300 -25 315 -10
rect 235 -50 275 -40
rect 235 -70 245 -50
rect 265 -70 275 -50
rect 235 -80 275 -70
<< polycont >>
rect 50 570 70 590
rect -55 385 -35 405
rect 60 350 80 370
rect 350 370 370 390
rect 180 180 200 200
rect 65 155 85 175
rect 350 200 370 220
rect 285 160 305 180
rect -35 -70 -15 -50
rect 245 -70 265 -50
<< locali >>
rect -45 710 -5 720
rect -45 640 -35 710
rect -15 640 -5 710
rect -45 630 -5 640
rect 60 710 150 720
rect 60 640 70 710
rect 90 640 120 710
rect 140 640 150 710
rect 60 630 150 640
rect 190 710 230 720
rect 190 640 200 710
rect 220 640 230 710
rect 190 630 230 640
rect 295 710 385 720
rect 295 640 305 710
rect 325 640 355 710
rect 375 640 385 710
rect 295 630 385 640
rect -45 610 -25 630
rect -85 590 -25 610
rect 40 590 80 600
rect 40 570 50 590
rect 70 570 80 590
rect 40 560 80 570
rect 40 530 60 560
rect 105 530 125 630
rect 315 610 335 630
rect 315 590 435 610
rect -45 520 -5 530
rect -45 450 -35 520
rect -15 450 -5 520
rect -45 440 -5 450
rect 20 520 60 530
rect 20 450 30 520
rect 50 450 60 520
rect 20 440 60 450
rect 85 520 125 530
rect 85 450 95 520
rect 115 450 125 520
rect 85 440 125 450
rect 190 520 230 530
rect 190 450 200 520
rect 220 450 230 520
rect 190 440 230 450
rect 295 520 335 530
rect 295 450 305 520
rect 325 450 335 520
rect 295 440 335 450
rect -45 415 -25 440
rect -65 405 -25 415
rect -65 385 -55 405
rect -35 385 -25 405
rect -65 375 -25 385
rect 40 400 60 440
rect 295 400 315 440
rect 40 380 70 400
rect 275 390 380 400
rect 275 380 350 390
rect 50 370 90 380
rect 50 350 60 370
rect 80 360 90 370
rect 80 350 140 360
rect 50 340 140 350
rect 275 340 295 380
rect 340 370 350 380
rect 370 370 380 390
rect 340 360 380 370
rect -45 310 -5 320
rect -45 240 -35 310
rect -15 240 -5 310
rect -45 230 -5 240
rect 60 310 100 320
rect 60 240 70 310
rect 90 240 100 310
rect 60 230 100 240
rect -45 210 -25 230
rect -65 190 -25 210
rect -65 85 -45 190
rect 75 185 95 230
rect 55 175 95 185
rect 55 155 65 175
rect 85 155 95 175
rect 55 145 95 155
rect 120 125 140 340
rect 190 330 230 340
rect 190 260 200 330
rect 220 260 230 330
rect 190 250 230 260
rect 255 330 295 340
rect 255 260 265 330
rect 285 260 295 330
rect 255 250 295 260
rect 320 330 360 340
rect 320 260 330 330
rect 350 260 360 330
rect 320 250 360 260
rect 190 210 210 250
rect 275 230 295 250
rect 275 220 380 230
rect 275 210 350 220
rect 170 200 210 210
rect 170 180 180 200
rect 200 180 210 200
rect 340 200 350 210
rect 370 200 380 220
rect 340 190 380 200
rect 170 170 210 180
rect 275 180 315 190
rect 275 160 285 180
rect 305 160 315 180
rect 275 150 315 160
rect 275 125 295 150
rect 400 125 420 590
rect 60 105 210 125
rect 60 85 80 105
rect 190 85 210 105
rect 275 105 420 125
rect 275 85 295 105
rect -65 75 -25 85
rect -65 5 -55 75
rect -35 5 -25 75
rect -65 -5 -25 5
rect 40 75 130 85
rect 40 5 50 75
rect 70 5 100 75
rect 120 5 130 75
rect 40 -5 130 5
rect 190 75 230 85
rect 190 5 200 75
rect 220 5 230 75
rect 190 -5 230 5
rect 255 75 295 85
rect 255 5 265 75
rect 285 5 295 75
rect 255 -5 295 5
rect 320 75 410 85
rect 320 5 330 75
rect 350 5 380 75
rect 400 5 410 75
rect 320 -5 410 5
rect -45 -50 -5 -40
rect -45 -70 -35 -50
rect -15 -70 -5 -50
rect -45 -80 -5 -70
rect 235 -50 275 -40
rect 235 -70 245 -50
rect 265 -70 275 -50
rect 235 -80 275 -70
<< viali >>
rect 70 640 90 710
rect 200 640 220 710
rect 95 450 115 520
rect 200 450 220 520
rect 330 260 350 330
rect 330 5 350 75
rect 380 5 400 75
rect -35 -70 -15 -50
rect 245 -70 265 -50
<< metal1 >>
rect -85 710 435 720
rect -85 640 70 710
rect 90 640 200 710
rect 220 640 435 710
rect -85 520 435 640
rect -85 450 95 520
rect 115 450 200 520
rect 220 450 435 520
rect -85 440 435 450
rect -85 330 435 340
rect -85 260 330 330
rect 350 260 435 330
rect -85 75 435 260
rect -85 5 330 75
rect 350 5 380 75
rect 400 5 435 75
rect -85 -10 435 5
rect -85 -50 435 -40
rect -85 -70 -35 -50
rect -15 -70 245 -50
rect 265 -70 435 -50
rect -85 -80 435 -70
<< labels >>
rlabel locali -85 600 -85 600 7 D
port 1 w
rlabel poly -85 390 -85 390 7 Db
port 2 w
rlabel metal1 -85 705 -85 705 7 VP
port 3 w
rlabel metal1 -85 15 -85 15 7 VN
port 4 w
rlabel metal1 -85 -60 -85 -60 7 clk
port 5 w
rlabel locali 435 600 435 600 3 Q
port 6 e
rlabel poly 435 390 435 390 3 Qb
port 7 e
<< end >>
