* SPICE3 file created from /home/madvlsi/Documents/Miniproject3/fcdiffamp_full.ext - technology: sky130A

.subckt fcdiffamp_layout V1 V2 VP VN Vcp Vbp Vcn Vbn Vout a_2400_2600#
X0 net5 Vcp net8 VP sky130_fd_pr__pfet_01v8 ad=7.5e+11p pd=6.5e+06u as=3e+12p ps=1.4e+07u w=3e+06u l=500000u
X1 a_400_0# V1 a_600_2600# VP sky130_fd_pr__pfet_01v8 ad=4.5e+12p pd=2.1e+07u as=1.05e+13p ps=4.9e+07u w=3e+06u l=500000u
X2 net8 Vcp net6 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X3 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=2.4e+13p pd=1.12e+08u as=0p ps=0u w=3e+06u l=500000u
X4 VP VP a_400_0# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X5 a_2400_2600# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=6e+12p pd=2.8e+07u as=1.2e+13p ps=5.6e+07u w=3e+06u l=500000u
X6 net6 net8 VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X7 Vout Vcp net11 VP sky130_fd_pr__pfet_01v8 ad=3e+12p pd=1.4e+07u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X8 a_2400_2600# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X9 a_400_0# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=6e+12p pd=2.8e+07u as=0p ps=0u w=3e+06u l=500000u
X10 VN Vbn a_400_0# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X11 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X12 net11 net8 VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X13 Vout VN VN VN sky130_fd_pr__nfet_01v8 ad=4.5e+12p pd=2.1e+07u as=0p ps=0u w=3e+06u l=500000u
X14 VP VP a_600_2600# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X15 Vout Vcn a_2400_2600# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X16 a_600_2600# V2 a_2400_2600# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3e+12p ps=1.4e+07u w=3e+06u l=500000u
X17 net8 Vcp net4 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X18 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X19 a_600_2600# Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X20 a_400_0# V1 a_600_2600# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X21 net4 net8 VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X22 VP net8 net5 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X23 VN VN net8 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.5e+12p ps=2.1e+07u w=3e+06u l=500000u
X24 a_2950_1200# Vcp Vout VP sky130_fd_pr__pfet_01v8 ad=7.5e+11p pd=6.5e+06u as=0p ps=0u w=3e+06u l=500000u
X25 net8 Vcn a_400_0# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X26 VP net8 a_1650_1200# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X27 VP net8 a_2950_1200# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X28 VN Vbn a_2400_2600# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X29 a_600_2600# Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X30 VN Vbn a_2400_2600# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X31 a_2400_2600# V2 a_600_2600# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X32 VN Vbn a_400_0# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X33 VP net8 net12 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X34 a_400_0# Vcn net8 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X35 VP Vbp a_600_2600# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X36 a_600_2600# V2 a_2400_2600# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X37 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X38 Vout Vcp a_2600_1200# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X39 a_400_0# VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X40 VP Vbp a_600_2600# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X41 Vout Vcn a_2400_2600# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X42 a_600_2600# V1 a_400_0# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X43 a_1650_1200# Vcp net8 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X44 a_2600_1200# net8 VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X45 net8 Vcn a_400_0# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X46 a_600_2600# V1 a_400_0# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X47 a_400_0# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X48 a_2400_2600# V2 a_600_2600# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X49 a_2400_2600# Vcn Vout VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X50 a_600_2600# VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X51 net12 Vcp Vout VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X52 a_2400_2600# Vcn Vout VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X53 a_400_0# Vcn net8 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X54 net8 VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X55 VN VN Vout VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
.ends

.subckt fc_bias VP VN Vbp Vbn Vcp Vcn
X0 net40 net39 net39 VN sky130_fd_pr__nfet_01v8 ad=1.95e+13p pd=9.1e+07u as=1.2e+13p ps=5.6e+07u w=3e+06u l=500000u
X1 a_900_3000# Vbp VP VP sky130_fd_pr__pfet_01v8 ad=1.5e+12p pd=7e+06u as=3.5265e+13p ps=1.681e+08u w=3e+06u l=500000u
X2 a_1700_0# Vbn a_n550_810# VN sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=6.5e+06u as=1.5e+12p ps=7e+06u w=3e+06u l=500000u
X3 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=2.985e+13p pd=1.399e+08u as=0p ps=0u w=3e+06u l=500000u
X4 Vbn Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3e+12p pd=1.4e+07u as=0p ps=0u w=3e+06u l=500000u
X5 net42 a_n550_810# a_n550_810# VP sky130_fd_pr__pfet_01v8 ad=1.8e+13p pd=8.4e+07u as=1.2e+13p ps=5.6e+07u w=3e+06u l=500000u
X6 net39 net39 net40 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X7 a_3650_0# Vbn a_3500_0# VN sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=6.5e+06u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X8 a_n550_810# a_n550_810# net42 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X9 Vbn Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3e+12p pd=1.4e+07u as=0p ps=0u w=3e+06u l=500000u
X10 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X11 VP Vbp net19 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X12 net40 net39 net39 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X13 net39 net39 net40 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X14 a_2450_3000# Vbp a_2300_3000# VP sky130_fd_pr__pfet_01v8 ad=7.5e+11p pd=6.5e+06u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X15 Vcp VP VP VP sky130_fd_pr__pfet_01v8 ad=4.5e+12p pd=2.1e+07u as=0p ps=0u w=3e+06u l=500000u
X16 VP Vbp Vcn VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3e+12p ps=1.4e+07u w=3e+06u l=500000u
X17 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X18 Vbp VP VP VP sky130_fd_pr__pfet_01v8 ad=3e+12p pd=1.4e+07u as=0p ps=0u w=3e+06u l=500000u
X19 a_4100_0# Vbn a_3950_0# VN sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=6.5e+06u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X20 net19 Vbp a_4250_3000# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X21 a_3800_0# Vbn a_3650_0# VN sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=6.5e+06u as=0p ps=0u w=3e+06u l=500000u
X22 VP VP Vcp VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X23 net40 Vcn Vcn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3e+12p ps=1.4e+07u w=3e+06u l=500000u
X24 a_n550_810# a_n550_810# net42 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X25 a_2300_3000# Vbp a_2150_3000# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X26 a_2750_0# Vbn a_2600_0# VN sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=6.5e+06u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X27 Vcp Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3e+12p pd=1.4e+07u as=0p ps=0u w=3e+06u l=500000u
X28 net42 a_n550_810# a_n550_810# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X29 a_2000_3000# Vbp a_1850_3000# VP sky130_fd_pr__pfet_01v8 ad=7.5e+11p pd=6.5e+06u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X30 net39 net39 net40 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X31 VP Vbp Vbp VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X32 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X33 a_n550_810# a_n550_810# net42 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X34 a_3200_0# Vbn a_3050_0# VN sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=6.5e+06u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X35 a_3350_3000# Vbp a_3200_3000# VP sky130_fd_pr__pfet_01v8 ad=7.5e+11p pd=6.5e+06u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X36 net40 net39 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X37 a_2900_0# Vbn a_2750_0# VN sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=6.5e+06u as=0p ps=0u w=3e+06u l=500000u
X38 a_2150_0# Vbn a_2000_0# VN sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=6.5e+06u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X39 net42 a_n550_810# a_n550_810# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X40 Vbn Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X41 a_3050_3000# Vbp a_2900_3000# VP sky130_fd_pr__pfet_01v8 ad=7.5e+11p pd=6.5e+06u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X42 a_1850_0# Vbn a_1700_0# VN sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=6.5e+06u as=0p ps=0u w=3e+06u l=500000u
X43 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X44 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X45 net39 net39 net40 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X46 net40 net39 net39 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X47 a_3200_3000# Vbp a_3050_3000# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X48 a_n550_810# VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X49 Vcn Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X50 VN Vbn Vbn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X51 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X52 VP VP a_900_3000# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X53 a_2900_3000# Vbp a_2750_3000# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X54 a_2300_0# Vbn a_2150_0# VN sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=6.5e+06u as=0p ps=0u w=3e+06u l=500000u
X55 Vcp Vcp net42 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X56 a_2000_0# Vbn a_1850_0# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X57 Vcn Vcn net40 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X58 net42 a_n550_810# VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X59 VP Vbp Vbn VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X60 a_4250_3000# Vbp a_4100_3000# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X61 net40 net39 net39 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X62 a_4250_0# Vbn a_4100_0# VN sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=6.5e+06u as=0p ps=0u w=3e+06u l=500000u
X63 a_n550_810# a_n550_810# net42 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X64 a_3950_0# Vbn a_3800_0# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X65 a_2150_3000# Vbp a_2000_3000# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X66 net40 net39 net39 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X67 Vbp Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X68 a_3950_3000# Vbp a_3800_3000# VP sky130_fd_pr__pfet_01v8 ad=7.5e+11p pd=6.5e+06u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X69 net39 net39 net40 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X70 net42 a_n550_810# VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X71 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X72 a_1850_3000# Vbp net1 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X73 a_4100_3000# Vbp a_3950_3000# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X74 VN net39 net40 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X75 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X76 net40 net39 net39 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X77 a_4400_0# Vbn a_4250_0# VN sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=6.5e+06u as=0p ps=0u w=3e+06u l=500000u
X78 a_n550_810# a_n550_810# net42 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X79 a_3800_3000# Vbp a_3650_3000# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X80 VN Vbn Vcp VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X81 net40 net39 net39 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X82 VP Vbp Vcn VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X83 Vcn Vcn net40 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X84 a_3350_0# Vbn a_3200_0# VN sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=6.5e+06u as=0p ps=0u w=3e+06u l=500000u
X85 net39 net39 net40 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X86 net1 Vbp net39 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.5e+12p ps=7e+06u w=3e+06u l=500000u
X87 a_3050_0# Vbn a_2900_0# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X88 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X89 VN Vbn Vbn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X90 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X91 VN net39 net40 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X92 a_n550_810# a_n550_810# net42 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X93 net42 Vcp Vcp VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X94 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X95 net40 Vcn Vcn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X96 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X97 net42 a_n550_810# a_n550_810# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X98 a_3500_0# Vbn a_3350_0# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X99 a_2750_3000# Vbp a_2600_3000# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X100 net39 net39 net40 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X101 net42 a_n550_810# a_n550_810# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X102 a_2450_0# Vbn a_2300_0# VN sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=6.5e+06u as=0p ps=0u w=3e+06u l=500000u
X103 a_n550_810# a_n550_810# net42 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X104 Vbn Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X105 VP Vbp Vbp VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X106 net40 net39 net39 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X107 VP a_n550_810# net42 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X108 a_2600_3000# Vbp a_2450_3000# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X109 net42 a_n550_810# a_n550_810# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X110 VP Vbp Vbn VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X111 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X112 net39 net39 net40 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X113 VN Vbn Vcp VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X114 net42 a_n550_810# a_n550_810# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X115 net42 Vcp Vcp VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X116 a_2600_0# Vbn a_2450_0# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X117 Vcn Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X118 net40 VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X119 net40 net39 VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X120 net39 VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X121 VP a_n550_810# net42 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X122 a_3650_3000# Vbp a_3500_3000# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.5e+11p ps=6.5e+06u w=3e+06u l=500000u
X123 VN Vbn a_4400_0# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X124 VN VN net40 VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X125 net42 a_n550_810# a_n550_810# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X126 Vcp Vcp net42 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X127 Vcp Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X128 a_n550_810# a_n550_810# net42 VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
X129 a_3500_3000# Vbp a_3350_3000# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=500000u
.ends

.subckt home/madvlsi/Documents/Miniproject3/fcdiffamp_full V1 V2 Vout Vcp Vcn Vbn
+ Vbp
Xfcdiffamp_layout_0 V1 V2 fc_bias_0/VP VSUBS Vcp Vbp Vcn Vbn Vout Vcp fcdiffamp_layout
Xfc_bias_0 fc_bias_0/VP VSUBS Vbp Vbn Vcp Vcn fc_bias
.ends

