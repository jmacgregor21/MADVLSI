magic
tech sky130A
timestamp 1614986124
<< nwell >>
rect -20 190 185 380
<< nmos >>
rect 50 0 65 100
<< pmos >>
rect 50 210 65 310
<< ndiff >>
rect 0 85 50 100
rect 0 15 15 85
rect 35 15 50 85
rect 0 0 50 15
rect 65 85 115 100
rect 65 15 80 85
rect 100 15 115 85
rect 65 0 115 15
<< pdiff >>
rect 0 295 50 310
rect 0 225 15 295
rect 35 225 50 295
rect 0 210 50 225
rect 65 295 115 310
rect 65 225 80 295
rect 100 225 115 295
rect 65 210 115 225
<< ndiffc >>
rect 15 15 35 85
rect 80 15 100 85
<< pdiffc >>
rect 15 225 35 295
rect 80 225 100 295
<< psubdiff >>
rect 115 85 165 100
rect 115 15 130 85
rect 150 15 165 85
rect 115 0 165 15
<< nsubdiff >>
rect 115 295 165 310
rect 115 225 130 295
rect 150 225 165 295
rect 115 210 165 225
<< psubdiffcont >>
rect 130 15 150 85
<< nsubdiffcont >>
rect 130 225 150 295
<< poly >>
rect 50 370 90 380
rect 50 350 60 370
rect 80 350 90 370
rect 50 340 90 350
rect 50 310 65 340
rect 50 100 65 210
rect 115 165 175 175
rect 115 145 125 165
rect 145 160 175 165
rect 145 145 155 160
rect 115 135 155 145
rect 50 -15 65 0
rect 0 -30 65 -15
<< polycont >>
rect 60 350 80 370
rect 125 145 145 165
<< locali >>
rect 50 370 185 380
rect 50 350 60 370
rect 80 360 185 370
rect 80 350 90 360
rect 50 340 90 350
rect 5 295 45 305
rect 5 225 15 295
rect 35 225 45 295
rect 5 215 45 225
rect 70 295 160 305
rect 70 225 80 295
rect 100 225 130 295
rect 150 225 160 295
rect 70 215 160 225
rect 5 155 25 215
rect 115 165 155 175
rect 115 155 125 165
rect 5 145 125 155
rect 145 145 155 165
rect 5 135 155 145
rect 5 95 25 135
rect 5 85 45 95
rect 5 15 15 85
rect 35 15 45 85
rect 5 5 45 15
rect 70 85 160 95
rect 70 15 80 85
rect 100 15 130 85
rect 150 15 160 85
rect 70 5 160 15
<< viali >>
rect 80 225 100 295
rect 130 225 150 295
rect 80 15 100 85
rect 130 15 150 85
<< metal1 >>
rect -20 295 185 340
rect -20 225 80 295
rect 100 225 130 295
rect 150 225 185 295
rect -20 205 185 225
rect 0 85 175 115
rect 0 15 80 85
rect 100 15 130 85
rect 150 15 175 85
rect 0 -35 175 15
<< labels >>
rlabel poly 0 -25 0 -25 7 A
port 1 w
rlabel poly 165 165 165 165 3 Y
port 2 e
rlabel metal1 0 -10 0 -10 7 VN
port 3 w
rlabel metal1 -20 235 -20 235 7 VP
port 4 w
<< end >>
