magic
tech sky130A
timestamp 1614543283
<< nwell >>
rect -145 645 465 825
rect -150 435 465 645
<< nmos >>
rect 0 245 15 345
rect 40 245 55 345
rect 105 245 120 345
rect 250 245 265 345
rect 315 245 330 345
rect 380 245 395 345
rect 0 0 15 100
rect 40 0 55 100
rect 105 0 120 100
rect 250 0 265 100
rect 315 0 330 100
rect 380 0 395 100
<< pmos >>
rect 0 705 15 805
rect 65 705 80 805
rect 130 705 145 805
rect 275 705 290 805
rect 315 705 330 805
rect 380 705 395 805
rect 0 460 15 560
rect 65 460 80 560
rect 130 460 145 560
rect 275 460 290 560
rect 315 460 330 560
rect 380 460 395 560
<< ndiff >>
rect -50 330 0 345
rect -50 260 -35 330
rect -15 260 0 330
rect -50 245 0 260
rect 15 245 40 345
rect 55 330 105 345
rect 55 260 70 330
rect 90 260 105 330
rect 55 245 105 260
rect 120 330 170 345
rect 120 260 135 330
rect 155 260 170 330
rect 120 245 170 260
rect 200 330 250 345
rect 200 260 215 330
rect 235 260 250 330
rect 200 245 250 260
rect 265 330 315 345
rect 265 260 280 330
rect 300 260 315 330
rect 265 245 315 260
rect 330 330 380 345
rect 330 260 345 330
rect 365 260 380 330
rect 330 245 380 260
rect 395 330 445 345
rect 395 260 410 330
rect 430 260 445 330
rect 395 245 445 260
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 0 40 100
rect 55 85 105 100
rect 55 15 70 85
rect 90 15 105 85
rect 55 0 105 15
rect 120 85 170 100
rect 120 15 135 85
rect 155 15 170 85
rect 120 0 170 15
rect 200 85 250 100
rect 200 15 215 85
rect 235 15 250 85
rect 200 0 250 15
rect 265 85 315 100
rect 265 15 280 85
rect 300 15 315 85
rect 265 0 315 15
rect 330 85 380 100
rect 330 15 345 85
rect 365 15 380 85
rect 330 0 380 15
rect 395 85 445 100
rect 395 15 410 85
rect 430 15 445 85
rect 395 0 445 15
<< pdiff >>
rect -50 790 0 805
rect -50 720 -35 790
rect -15 720 0 790
rect -50 705 0 720
rect 15 790 65 805
rect 15 720 30 790
rect 50 720 65 790
rect 15 705 65 720
rect 80 790 130 805
rect 80 720 95 790
rect 115 720 130 790
rect 80 705 130 720
rect 145 790 195 805
rect 145 720 160 790
rect 180 720 195 790
rect 145 705 195 720
rect 225 790 275 805
rect 225 720 240 790
rect 260 720 275 790
rect 225 705 275 720
rect 290 705 315 805
rect 330 790 380 805
rect 330 720 345 790
rect 365 720 380 790
rect 330 705 380 720
rect 395 790 445 805
rect 395 720 410 790
rect 430 720 445 790
rect 395 705 445 720
rect -50 545 0 560
rect -50 475 -35 545
rect -15 475 0 545
rect -50 460 0 475
rect 15 545 65 560
rect 15 475 30 545
rect 50 475 65 545
rect 15 460 65 475
rect 80 545 130 560
rect 80 475 95 545
rect 115 475 130 545
rect 80 460 130 475
rect 145 545 195 560
rect 145 475 160 545
rect 180 475 195 545
rect 145 460 195 475
rect 225 545 275 560
rect 225 475 240 545
rect 260 475 275 545
rect 225 460 275 475
rect 290 460 315 560
rect 330 545 380 560
rect 330 475 345 545
rect 365 475 380 545
rect 330 460 380 475
rect 395 545 445 560
rect 395 475 410 545
rect 430 475 445 545
rect 395 460 445 475
<< ndiffc >>
rect -35 260 -15 330
rect 70 260 90 330
rect 135 260 155 330
rect 215 260 235 330
rect 280 260 300 330
rect 345 260 365 330
rect 410 260 430 330
rect -35 15 -15 85
rect 70 15 90 85
rect 135 15 155 85
rect 215 15 235 85
rect 280 15 300 85
rect 345 15 365 85
rect 410 15 430 85
<< pdiffc >>
rect -35 720 -15 790
rect 30 720 50 790
rect 95 720 115 790
rect 160 720 180 790
rect 240 720 260 790
rect 345 720 365 790
rect 410 720 430 790
rect -35 475 -15 545
rect 30 475 50 545
rect 95 475 115 545
rect 160 475 180 545
rect 240 475 260 545
rect 345 475 365 545
rect 410 475 430 545
<< psubdiff >>
rect -130 85 -80 100
rect -130 15 -115 85
rect -95 15 -80 85
rect -130 0 -80 15
<< nsubdiff >>
rect -130 545 -80 560
rect -130 475 -115 545
rect -95 475 -80 545
rect -130 460 -80 475
<< psubdiffcont >>
rect -115 15 -95 85
<< nsubdiffcont >>
rect -115 475 -95 545
<< poly >>
rect 0 805 15 820
rect 65 805 80 820
rect 130 805 145 820
rect 275 805 290 820
rect 315 805 330 820
rect 380 805 395 820
rect 0 695 15 705
rect -50 680 15 695
rect 0 560 15 575
rect 65 560 80 705
rect 130 690 145 705
rect 275 690 290 705
rect 105 680 145 690
rect 105 660 115 680
rect 135 660 145 680
rect 105 650 145 660
rect 170 680 290 690
rect 170 660 180 680
rect 200 675 290 680
rect 200 660 210 675
rect 170 650 210 660
rect 170 590 185 650
rect 130 575 185 590
rect 130 560 145 575
rect 275 560 290 575
rect 315 560 330 705
rect 380 690 395 705
rect 420 680 465 695
rect 420 615 435 680
rect 355 605 435 615
rect 355 585 365 605
rect 385 600 435 605
rect 385 585 395 600
rect 355 575 395 585
rect 380 560 395 575
rect 0 400 15 460
rect 65 450 80 460
rect -25 390 15 400
rect -25 370 -15 390
rect 5 370 15 390
rect -25 360 15 370
rect 0 345 15 360
rect 40 435 80 450
rect 130 445 145 460
rect 275 445 290 460
rect 40 345 55 435
rect 105 430 145 445
rect 250 435 290 445
rect 105 345 120 430
rect 250 415 260 435
rect 280 415 290 435
rect 250 405 290 415
rect 250 345 265 405
rect 315 345 330 460
rect 380 345 395 460
rect 0 230 15 245
rect -50 110 15 125
rect 0 100 15 110
rect 40 100 55 245
rect 105 230 120 245
rect 250 230 265 245
rect 80 220 120 230
rect 80 200 90 220
rect 110 205 120 220
rect 110 200 160 205
rect 80 190 160 200
rect 145 130 160 190
rect 145 115 265 130
rect 105 100 120 115
rect 250 100 265 115
rect 315 100 330 245
rect 380 230 395 245
rect 380 215 435 230
rect 355 145 395 155
rect 355 125 365 145
rect 385 125 395 145
rect 355 115 395 125
rect 380 100 395 115
rect 420 150 435 215
rect 420 140 460 150
rect 420 120 430 140
rect 450 120 460 140
rect 420 110 460 120
rect 0 -15 15 0
rect 40 -15 55 0
rect 105 -15 120 0
rect 250 -15 265 0
rect 315 -15 330 0
rect 380 -15 395 0
rect 80 -25 120 -15
rect 80 -45 90 -25
rect 110 -45 120 -25
rect 80 -55 120 -45
<< polycont >>
rect 115 660 135 680
rect 180 660 200 680
rect 365 585 385 605
rect -15 370 5 390
rect 260 415 280 435
rect 90 200 110 220
rect 365 125 385 145
rect 430 120 450 140
rect 90 -45 110 -25
<< locali >>
rect -25 820 105 840
rect -25 800 -5 820
rect 85 800 105 820
rect -45 790 -5 800
rect -45 720 -35 790
rect -15 720 -5 790
rect -45 710 -5 720
rect 20 790 60 800
rect 20 720 30 790
rect 50 720 60 790
rect 20 710 60 720
rect 85 790 125 800
rect 85 720 95 790
rect 115 720 125 790
rect 85 710 125 720
rect 150 790 190 800
rect 150 720 160 790
rect 180 720 190 790
rect 150 710 190 720
rect 230 790 270 800
rect 230 720 240 790
rect 260 720 270 790
rect 230 710 270 720
rect 335 790 375 800
rect 335 720 345 790
rect 365 720 375 790
rect 335 710 375 720
rect 400 790 440 800
rect 400 720 410 790
rect 430 720 440 790
rect 400 710 440 720
rect 20 555 40 710
rect 170 690 190 710
rect 105 680 145 690
rect 105 660 115 680
rect 135 660 145 680
rect 105 650 145 660
rect 170 680 210 690
rect 170 660 180 680
rect 200 660 210 680
rect 170 650 210 660
rect 125 595 145 650
rect 355 615 375 710
rect 355 605 395 615
rect 125 575 170 595
rect 355 585 365 605
rect 385 585 395 605
rect 355 575 395 585
rect 150 555 170 575
rect 420 555 440 710
rect -125 545 -85 555
rect -125 475 -115 545
rect -95 475 -85 545
rect -125 465 -85 475
rect -45 545 -5 555
rect -45 475 -35 545
rect -15 475 -5 545
rect -45 465 -5 475
rect 20 545 60 555
rect 20 475 30 545
rect 50 475 60 545
rect 20 465 60 475
rect 85 545 125 555
rect 85 475 95 545
rect 115 475 125 545
rect 85 465 125 475
rect 150 545 190 555
rect 150 475 160 545
rect 180 475 190 545
rect 150 465 190 475
rect 230 545 270 555
rect 230 475 240 545
rect 260 475 270 545
rect 230 465 270 475
rect 335 545 375 555
rect 335 475 345 545
rect 365 475 375 545
rect 335 465 375 475
rect 400 545 440 555
rect 400 475 410 545
rect 430 475 440 545
rect 400 465 440 475
rect -25 445 -5 465
rect 85 445 105 465
rect -25 425 105 445
rect 150 445 170 465
rect 355 445 375 465
rect 150 435 290 445
rect 150 425 260 435
rect -25 390 15 400
rect -25 380 -15 390
rect -45 370 -15 380
rect 5 370 15 390
rect 150 380 170 425
rect 250 415 260 425
rect 280 415 290 435
rect 355 425 440 445
rect 250 405 290 415
rect 420 380 440 425
rect -45 360 15 370
rect 80 360 170 380
rect 225 360 355 380
rect 80 340 100 360
rect 225 340 245 360
rect 335 340 355 360
rect 420 360 465 380
rect 420 340 440 360
rect -45 330 -5 340
rect -45 260 -35 330
rect -15 260 -5 330
rect 60 330 100 340
rect 60 270 70 330
rect -45 250 -5 260
rect 20 260 70 270
rect 90 260 100 330
rect 20 250 100 260
rect 125 330 165 340
rect 125 260 135 330
rect 155 260 165 330
rect 125 250 165 260
rect 205 330 245 340
rect 205 260 215 330
rect 235 260 245 330
rect 205 250 245 260
rect 270 330 310 340
rect 270 260 280 330
rect 300 260 310 330
rect 270 250 310 260
rect 335 330 375 340
rect 335 260 345 330
rect 365 260 375 330
rect 335 250 375 260
rect 400 330 440 340
rect 400 260 410 330
rect 430 260 440 330
rect 400 250 440 260
rect -45 95 -25 250
rect -125 85 -85 95
rect -125 15 -115 85
rect -95 15 -85 85
rect -125 5 -85 15
rect -45 85 -5 95
rect -45 15 -35 85
rect -15 15 -5 85
rect -45 5 -5 15
rect 20 -15 40 250
rect 80 220 120 230
rect 80 200 90 220
rect 110 200 120 220
rect 80 190 120 200
rect 80 95 100 190
rect 145 95 165 250
rect 270 95 295 250
rect 400 230 420 250
rect 375 210 420 230
rect 375 155 395 210
rect 355 145 395 155
rect 355 125 365 145
rect 385 125 395 145
rect 355 115 395 125
rect 420 140 460 150
rect 420 120 430 140
rect 450 120 460 140
rect 420 110 460 120
rect 420 95 440 110
rect 60 85 100 95
rect 60 15 70 85
rect 90 15 100 85
rect 60 5 100 15
rect 125 85 165 95
rect 125 15 135 85
rect 155 15 165 85
rect 125 5 165 15
rect 205 85 245 95
rect 205 15 215 85
rect 235 15 245 85
rect 205 5 245 15
rect 270 85 310 95
rect 270 15 280 85
rect 300 15 310 85
rect 270 5 310 15
rect 335 85 375 95
rect 335 15 345 85
rect 365 15 375 85
rect 335 5 375 15
rect 400 85 440 95
rect 400 15 410 85
rect 430 15 440 85
rect 400 5 440 15
rect 225 -15 245 5
rect 335 -15 355 5
rect 20 -25 120 -15
rect 20 -35 90 -25
rect 80 -45 90 -35
rect 110 -45 120 -25
rect 225 -35 355 -15
rect 80 -55 120 -45
<< end >>
