magic
tech sky130A
timestamp 1615160756
<< nwell >>
rect -60 975 2235 1165
rect -60 475 2235 815
<< nmos >>
rect 65 -5 115 295
rect 165 -5 215 295
rect 265 -5 315 295
rect 365 -5 415 295
rect 465 -5 515 295
rect 565 -5 615 295
rect 665 -5 715 295
rect 765 -5 815 295
rect 865 -5 915 295
rect 965 -5 1015 295
rect 1165 -5 1215 295
rect 1265 -5 1315 295
rect 1365 -5 1415 295
rect 1465 -5 1515 295
rect 1565 -5 1615 295
rect 1665 -5 1715 295
rect 1765 -5 1815 295
rect 1865 -5 1915 295
rect 1965 -5 2015 295
rect 2065 -5 2115 295
<< pmos >>
rect 65 995 115 1145
rect 165 995 215 1145
rect 265 995 315 1145
rect 365 995 415 1145
rect 465 995 515 1145
rect 565 995 615 1145
rect 665 995 715 1145
rect 765 995 815 1145
rect 865 995 915 1145
rect 965 995 1015 1145
rect 1165 995 1215 1145
rect 1265 995 1315 1145
rect 1365 995 1415 1145
rect 1465 995 1515 1145
rect 1565 995 1615 1145
rect 1665 995 1715 1145
rect 1765 995 1815 1145
rect 1865 995 1915 1145
rect 1965 995 2015 1145
rect 2065 995 2115 1145
rect 65 495 115 795
rect 165 495 215 795
rect 265 495 315 795
rect 365 495 415 795
rect 465 495 515 795
rect 565 495 615 795
rect 665 495 715 795
rect 765 495 815 795
rect 865 495 915 795
rect 965 495 1015 795
rect 1165 495 1215 795
rect 1265 495 1315 795
rect 1365 495 1415 795
rect 1465 495 1515 795
rect 1565 495 1615 795
rect 1665 495 1715 795
rect 1765 495 1815 795
rect 1865 495 1915 795
rect 1965 495 2015 795
rect 2065 495 2115 795
<< ndiff >>
rect 15 280 65 295
rect 15 10 30 280
rect 50 10 65 280
rect 15 -5 65 10
rect 115 280 165 295
rect 115 10 130 280
rect 150 10 165 280
rect 115 -5 165 10
rect 215 280 265 295
rect 215 10 230 280
rect 250 10 265 280
rect 215 -5 265 10
rect 315 280 365 295
rect 315 10 330 280
rect 350 10 365 280
rect 315 -5 365 10
rect 415 280 465 295
rect 415 10 430 280
rect 450 10 465 280
rect 415 -5 465 10
rect 515 280 565 295
rect 515 10 530 280
rect 550 10 565 280
rect 515 -5 565 10
rect 615 280 665 295
rect 615 10 630 280
rect 650 10 665 280
rect 615 -5 665 10
rect 715 280 765 295
rect 715 10 730 280
rect 750 10 765 280
rect 715 -5 765 10
rect 815 280 865 295
rect 815 10 830 280
rect 850 10 865 280
rect 815 -5 865 10
rect 915 280 965 295
rect 915 10 930 280
rect 950 10 965 280
rect 915 -5 965 10
rect 1015 280 1065 295
rect 1115 280 1165 295
rect 1015 10 1030 280
rect 1050 10 1065 280
rect 1115 10 1130 280
rect 1150 10 1165 280
rect 1015 -5 1065 10
rect 1115 -5 1165 10
rect 1215 280 1265 295
rect 1215 10 1230 280
rect 1250 10 1265 280
rect 1215 -5 1265 10
rect 1315 280 1365 295
rect 1315 10 1330 280
rect 1350 10 1365 280
rect 1315 -5 1365 10
rect 1415 280 1465 295
rect 1415 10 1430 280
rect 1450 10 1465 280
rect 1415 -5 1465 10
rect 1515 280 1565 295
rect 1515 10 1530 280
rect 1550 10 1565 280
rect 1515 -5 1565 10
rect 1615 280 1665 295
rect 1615 10 1630 280
rect 1650 10 1665 280
rect 1615 -5 1665 10
rect 1715 280 1765 295
rect 1715 10 1730 280
rect 1750 10 1765 280
rect 1715 -5 1765 10
rect 1815 280 1865 295
rect 1815 10 1830 280
rect 1850 10 1865 280
rect 1815 -5 1865 10
rect 1915 280 1965 295
rect 1915 10 1930 280
rect 1950 10 1965 280
rect 1915 -5 1965 10
rect 2015 280 2065 295
rect 2015 10 2030 280
rect 2050 10 2065 280
rect 2015 -5 2065 10
rect 2115 280 2165 295
rect 2115 10 2130 280
rect 2150 10 2165 280
rect 2115 -5 2165 10
<< pdiff >>
rect 15 1130 65 1145
rect 15 1010 30 1130
rect 50 1010 65 1130
rect 15 995 65 1010
rect 115 1130 165 1145
rect 115 1010 130 1130
rect 150 1010 165 1130
rect 115 995 165 1010
rect 215 1130 265 1145
rect 215 1010 230 1130
rect 250 1010 265 1130
rect 215 995 265 1010
rect 315 1130 365 1145
rect 315 1010 330 1130
rect 350 1010 365 1130
rect 315 995 365 1010
rect 415 1130 465 1145
rect 415 1010 430 1130
rect 450 1010 465 1130
rect 415 995 465 1010
rect 515 1130 565 1145
rect 515 1010 530 1130
rect 550 1010 565 1130
rect 515 995 565 1010
rect 615 1130 665 1145
rect 615 1010 630 1130
rect 650 1010 665 1130
rect 615 995 665 1010
rect 715 1130 765 1145
rect 715 1010 730 1130
rect 750 1010 765 1130
rect 715 995 765 1010
rect 815 1130 865 1145
rect 815 1010 830 1130
rect 850 1010 865 1130
rect 815 995 865 1010
rect 915 1130 965 1145
rect 915 1010 930 1130
rect 950 1010 965 1130
rect 915 995 965 1010
rect 1015 1130 1065 1145
rect 1115 1130 1165 1145
rect 1015 1010 1030 1130
rect 1050 1010 1065 1130
rect 1115 1010 1130 1130
rect 1150 1010 1165 1130
rect 1015 995 1065 1010
rect 1115 995 1165 1010
rect 1215 1130 1265 1145
rect 1215 1010 1230 1130
rect 1250 1010 1265 1130
rect 1215 995 1265 1010
rect 1315 1130 1365 1145
rect 1315 1010 1330 1130
rect 1350 1010 1365 1130
rect 1315 995 1365 1010
rect 1415 1130 1465 1145
rect 1415 1010 1430 1130
rect 1450 1010 1465 1130
rect 1415 995 1465 1010
rect 1515 1130 1565 1145
rect 1515 1010 1530 1130
rect 1550 1010 1565 1130
rect 1515 995 1565 1010
rect 1615 1130 1665 1145
rect 1615 1010 1630 1130
rect 1650 1010 1665 1130
rect 1615 995 1665 1010
rect 1715 1130 1765 1145
rect 1715 1010 1730 1130
rect 1750 1010 1765 1130
rect 1715 995 1765 1010
rect 1815 1130 1865 1145
rect 1815 1010 1830 1130
rect 1850 1010 1865 1130
rect 1815 995 1865 1010
rect 1915 1130 1965 1145
rect 1915 1010 1930 1130
rect 1950 1010 1965 1130
rect 1915 995 1965 1010
rect 2015 1130 2065 1145
rect 2015 1010 2030 1130
rect 2050 1010 2065 1130
rect 2015 995 2065 1010
rect 2115 1130 2165 1145
rect 2115 1010 2130 1130
rect 2150 1010 2165 1130
rect 2115 995 2165 1010
rect 15 780 65 795
rect 15 510 30 780
rect 50 510 65 780
rect 15 495 65 510
rect 115 780 165 795
rect 115 510 130 780
rect 150 510 165 780
rect 115 495 165 510
rect 215 780 265 795
rect 215 510 230 780
rect 250 510 265 780
rect 215 495 265 510
rect 315 780 365 795
rect 315 510 330 780
rect 350 510 365 780
rect 315 495 365 510
rect 415 780 465 795
rect 415 510 430 780
rect 450 510 465 780
rect 415 495 465 510
rect 515 780 565 795
rect 515 510 530 780
rect 550 510 565 780
rect 515 495 565 510
rect 615 780 665 795
rect 615 510 630 780
rect 650 510 665 780
rect 615 495 665 510
rect 715 780 765 795
rect 715 510 730 780
rect 750 510 765 780
rect 715 495 765 510
rect 815 780 865 795
rect 815 510 830 780
rect 850 510 865 780
rect 815 495 865 510
rect 915 780 965 795
rect 915 510 930 780
rect 950 510 965 780
rect 915 495 965 510
rect 1015 780 1065 795
rect 1115 780 1165 795
rect 1015 510 1030 780
rect 1050 510 1065 780
rect 1115 510 1130 780
rect 1150 510 1165 780
rect 1015 495 1065 510
rect 1115 495 1165 510
rect 1215 780 1265 795
rect 1215 510 1230 780
rect 1250 510 1265 780
rect 1215 495 1265 510
rect 1315 780 1365 795
rect 1315 510 1330 780
rect 1350 510 1365 780
rect 1315 495 1365 510
rect 1415 780 1465 795
rect 1415 510 1430 780
rect 1450 510 1465 780
rect 1415 495 1465 510
rect 1515 780 1565 795
rect 1515 510 1530 780
rect 1550 510 1565 780
rect 1515 495 1565 510
rect 1615 780 1665 795
rect 1615 510 1630 780
rect 1650 510 1665 780
rect 1615 495 1665 510
rect 1715 780 1765 795
rect 1715 510 1730 780
rect 1750 510 1765 780
rect 1715 495 1765 510
rect 1815 780 1865 795
rect 1815 510 1830 780
rect 1850 510 1865 780
rect 1815 495 1865 510
rect 1915 780 1965 795
rect 1915 510 1930 780
rect 1950 510 1965 780
rect 1915 495 1965 510
rect 2015 780 2065 795
rect 2015 510 2030 780
rect 2050 510 2065 780
rect 2015 495 2065 510
rect 2115 780 2165 795
rect 2115 510 2130 780
rect 2150 510 2165 780
rect 2115 495 2165 510
<< ndiffc >>
rect 30 10 50 280
rect 130 10 150 280
rect 230 10 250 280
rect 330 10 350 280
rect 430 10 450 280
rect 530 10 550 280
rect 630 10 650 280
rect 730 10 750 280
rect 830 10 850 280
rect 930 10 950 280
rect 1030 10 1050 280
rect 1130 10 1150 280
rect 1230 10 1250 280
rect 1330 10 1350 280
rect 1430 10 1450 280
rect 1530 10 1550 280
rect 1630 10 1650 280
rect 1730 10 1750 280
rect 1830 10 1850 280
rect 1930 10 1950 280
rect 2030 10 2050 280
rect 2130 10 2150 280
<< pdiffc >>
rect 30 1010 50 1130
rect 130 1010 150 1130
rect 230 1010 250 1130
rect 330 1010 350 1130
rect 430 1010 450 1130
rect 530 1010 550 1130
rect 630 1010 650 1130
rect 730 1010 750 1130
rect 830 1010 850 1130
rect 930 1010 950 1130
rect 1030 1010 1050 1130
rect 1130 1010 1150 1130
rect 1230 1010 1250 1130
rect 1330 1010 1350 1130
rect 1430 1010 1450 1130
rect 1530 1010 1550 1130
rect 1630 1010 1650 1130
rect 1730 1010 1750 1130
rect 1830 1010 1850 1130
rect 1930 1010 1950 1130
rect 2030 1010 2050 1130
rect 2130 1010 2150 1130
rect 30 510 50 780
rect 130 510 150 780
rect 230 510 250 780
rect 330 510 350 780
rect 430 510 450 780
rect 530 510 550 780
rect 630 510 650 780
rect 730 510 750 780
rect 830 510 850 780
rect 930 510 950 780
rect 1030 510 1050 780
rect 1130 510 1150 780
rect 1230 510 1250 780
rect 1330 510 1350 780
rect 1430 510 1450 780
rect 1530 510 1550 780
rect 1630 510 1650 780
rect 1730 510 1750 780
rect 1830 510 1850 780
rect 1930 510 1950 780
rect 2030 510 2050 780
rect 2130 510 2150 780
<< psubdiff >>
rect -40 280 15 295
rect -40 10 -25 280
rect 0 10 15 280
rect -40 -5 15 10
rect 1065 280 1115 295
rect 1065 10 1080 280
rect 1100 10 1115 280
rect 1065 -5 1115 10
rect 2165 280 2215 295
rect 2165 10 2180 280
rect 2200 10 2215 280
rect 2165 -5 2215 10
<< nsubdiff >>
rect -40 1130 15 1145
rect -40 1010 -25 1130
rect 0 1010 15 1130
rect -40 995 15 1010
rect 1065 1130 1115 1145
rect 1065 1010 1080 1130
rect 1100 1010 1115 1130
rect 1065 995 1115 1010
rect 2165 1130 2215 1145
rect 2165 1010 2180 1130
rect 2200 1010 2215 1130
rect 2165 995 2215 1010
rect -40 780 15 795
rect -40 510 -25 780
rect 0 510 15 780
rect -40 495 15 510
rect 1065 780 1115 795
rect 1065 510 1080 780
rect 1100 510 1115 780
rect 1065 495 1115 510
rect 2165 780 2215 795
rect 2165 510 2180 780
rect 2200 510 2215 780
rect 2165 495 2215 510
<< psubdiffcont >>
rect -25 10 0 280
rect 1080 10 1100 280
rect 2180 10 2200 280
<< nsubdiffcont >>
rect -25 1010 0 1130
rect 1080 1010 1100 1130
rect 2180 1010 2200 1130
rect -25 510 0 780
rect 1080 510 1100 780
rect 2180 510 2200 780
<< poly >>
rect 165 1190 215 1205
rect 165 1170 180 1190
rect 200 1170 215 1190
rect 65 1145 115 1160
rect 165 1145 215 1170
rect 265 1190 315 1205
rect 265 1170 280 1190
rect 300 1170 315 1190
rect 265 1145 315 1170
rect 365 1190 415 1205
rect 365 1170 380 1190
rect 400 1170 415 1190
rect 365 1145 415 1170
rect 465 1190 515 1205
rect 465 1170 480 1190
rect 500 1170 515 1190
rect 465 1145 515 1170
rect 565 1190 615 1205
rect 565 1170 580 1190
rect 600 1170 615 1190
rect 565 1145 615 1170
rect 665 1190 715 1205
rect 665 1170 680 1190
rect 700 1170 715 1190
rect 665 1145 715 1170
rect 765 1190 815 1205
rect 765 1170 780 1190
rect 800 1170 815 1190
rect 765 1145 815 1170
rect 865 1190 915 1205
rect 865 1170 880 1190
rect 900 1170 915 1190
rect 865 1145 915 1170
rect 1265 1190 1315 1205
rect 1265 1170 1280 1190
rect 1300 1170 1315 1190
rect 965 1145 1015 1160
rect 1165 1145 1215 1160
rect 1265 1145 1315 1170
rect 1365 1190 1415 1205
rect 1365 1170 1380 1190
rect 1400 1170 1415 1190
rect 1365 1145 1415 1170
rect 1465 1190 1515 1205
rect 1465 1170 1480 1190
rect 1500 1170 1515 1190
rect 1465 1145 1515 1170
rect 1565 1190 1615 1205
rect 1565 1170 1580 1190
rect 1600 1170 1615 1190
rect 1565 1145 1615 1170
rect 1665 1190 1715 1205
rect 1665 1170 1680 1190
rect 1700 1170 1715 1190
rect 1665 1145 1715 1170
rect 1765 1190 1815 1205
rect 1765 1170 1780 1190
rect 1800 1170 1815 1190
rect 1765 1145 1815 1170
rect 1865 1190 1915 1205
rect 1865 1170 1880 1190
rect 1900 1170 1915 1190
rect 1865 1145 1915 1170
rect 1965 1190 2015 1205
rect 1965 1170 1980 1190
rect 2000 1170 2015 1190
rect 1965 1145 2015 1170
rect 2065 1145 2115 1160
rect 65 985 115 995
rect 20 970 115 985
rect 165 980 215 995
rect 265 980 315 995
rect 365 980 415 995
rect 465 980 515 995
rect 565 980 615 995
rect 665 980 715 995
rect 765 980 815 995
rect 865 980 915 995
rect 965 985 1015 995
rect 1165 985 1215 995
rect 965 970 1215 985
rect 1265 980 1315 995
rect 1365 980 1415 995
rect 1465 980 1515 995
rect 1565 980 1615 995
rect 1665 980 1715 995
rect 1765 980 1815 995
rect 1865 980 1915 995
rect 1965 980 2015 995
rect 2065 985 2115 995
rect 2065 970 2160 985
rect 20 950 30 970
rect 50 950 60 970
rect 20 940 60 950
rect 1070 950 1080 970
rect 1100 950 1110 970
rect 1070 940 1110 950
rect 2120 950 2130 970
rect 2150 950 2160 970
rect 2120 940 2160 950
rect 20 840 60 850
rect 20 820 30 840
rect 50 820 60 840
rect 1070 840 1110 850
rect 1070 820 1080 840
rect 1100 820 1110 840
rect 1265 840 1315 855
rect 1265 820 1280 840
rect 1300 820 1315 840
rect 20 805 115 820
rect 65 795 115 805
rect 165 795 215 810
rect 265 795 315 810
rect 365 795 415 810
rect 465 795 515 810
rect 565 795 615 810
rect 665 795 715 810
rect 765 795 815 810
rect 865 795 915 810
rect 965 805 1215 820
rect 965 795 1015 805
rect 1165 795 1215 805
rect 1265 795 1315 820
rect 1365 840 1415 855
rect 1365 820 1380 840
rect 1400 820 1415 840
rect 1365 795 1415 820
rect 1465 840 1515 855
rect 1465 820 1480 840
rect 1500 820 1515 840
rect 1465 795 1515 820
rect 1565 840 1615 855
rect 1565 820 1580 840
rect 1600 820 1615 840
rect 1565 795 1615 820
rect 1665 840 1715 855
rect 1665 820 1680 840
rect 1700 820 1715 840
rect 1665 795 1715 820
rect 1765 840 1815 855
rect 1765 820 1780 840
rect 1800 820 1815 840
rect 1765 795 1815 820
rect 1865 840 1915 855
rect 1865 820 1880 840
rect 1900 820 1915 840
rect 1865 795 1915 820
rect 1965 840 2015 855
rect 1965 820 1980 840
rect 2000 820 2015 840
rect 2120 840 2160 850
rect 2120 820 2130 840
rect 2150 820 2160 840
rect 1965 795 2015 820
rect 2065 805 2160 820
rect 2065 795 2115 805
rect 65 480 115 495
rect 165 480 215 495
rect 265 480 315 495
rect 365 480 415 495
rect 465 480 515 495
rect 565 480 615 495
rect 665 480 715 495
rect 765 480 815 495
rect 865 480 915 495
rect 965 480 1015 495
rect 1165 480 1215 495
rect 1265 480 1315 495
rect 1365 480 1415 495
rect 1465 480 1515 495
rect 1565 480 1615 495
rect 1665 480 1715 495
rect 1765 480 1815 495
rect 1865 480 1915 495
rect 1965 480 2015 495
rect 2065 480 2115 495
rect 65 295 115 310
rect 165 295 215 310
rect 265 295 315 310
rect 365 295 415 310
rect 465 295 515 310
rect 565 295 615 310
rect 665 295 715 310
rect 765 295 815 310
rect 865 295 915 310
rect 965 295 1015 310
rect 1165 295 1215 310
rect 1265 295 1315 310
rect 1365 295 1415 310
rect 1465 295 1515 310
rect 1565 295 1615 310
rect 1665 295 1715 310
rect 1765 295 1815 310
rect 1865 295 1915 310
rect 1965 295 2015 310
rect 2065 295 2115 310
rect 65 -15 115 -5
rect 20 -30 115 -15
rect 20 -35 60 -30
rect 20 -55 30 -35
rect 50 -55 60 -35
rect 20 -65 60 -55
rect 165 -35 215 -5
rect 165 -55 180 -35
rect 200 -55 215 -35
rect 165 -70 215 -55
rect 265 -35 315 -5
rect 265 -55 280 -35
rect 300 -55 315 -35
rect 265 -70 315 -55
rect 365 -35 415 -5
rect 365 -55 380 -35
rect 400 -55 415 -35
rect 365 -70 415 -55
rect 465 -35 515 -5
rect 465 -55 480 -35
rect 500 -55 515 -35
rect 465 -70 515 -55
rect 565 -35 615 -5
rect 565 -55 580 -35
rect 600 -55 615 -35
rect 565 -70 615 -55
rect 665 -35 715 -5
rect 665 -55 680 -35
rect 700 -55 715 -35
rect 665 -70 715 -55
rect 765 -35 815 -5
rect 765 -55 780 -35
rect 800 -55 815 -35
rect 765 -70 815 -55
rect 865 -35 915 -5
rect 965 -15 1015 -5
rect 1165 -15 1215 -5
rect 965 -30 1215 -15
rect 1265 -30 1315 -5
rect 865 -55 880 -35
rect 900 -55 915 -35
rect 865 -70 915 -55
rect 1070 -50 1080 -30
rect 1100 -50 1110 -30
rect 1070 -60 1110 -50
rect 1265 -50 1280 -30
rect 1300 -50 1315 -30
rect 1265 -65 1315 -50
rect 1365 -30 1415 -5
rect 1365 -50 1380 -30
rect 1400 -50 1415 -30
rect 1365 -65 1415 -50
rect 1465 -30 1515 -5
rect 1465 -50 1480 -30
rect 1500 -50 1515 -30
rect 1465 -65 1515 -50
rect 1565 -30 1615 -5
rect 1565 -50 1580 -30
rect 1600 -50 1615 -30
rect 1565 -65 1615 -50
rect 1665 -30 1715 -5
rect 1665 -50 1680 -30
rect 1700 -50 1715 -30
rect 1665 -65 1715 -50
rect 1765 -30 1815 -5
rect 1765 -50 1780 -30
rect 1800 -50 1815 -30
rect 1765 -65 1815 -50
rect 1865 -30 1915 -5
rect 1865 -50 1880 -30
rect 1900 -50 1915 -30
rect 1865 -65 1915 -50
rect 1965 -30 2015 -5
rect 2065 -15 2115 -5
rect 2065 -30 2160 -15
rect 1965 -50 1980 -30
rect 2000 -50 2015 -30
rect 1965 -65 2015 -50
rect 2120 -50 2130 -30
rect 2150 -50 2160 -30
rect 2120 -60 2160 -50
<< polycont >>
rect 180 1170 200 1190
rect 280 1170 300 1190
rect 380 1170 400 1190
rect 480 1170 500 1190
rect 580 1170 600 1190
rect 680 1170 700 1190
rect 780 1170 800 1190
rect 880 1170 900 1190
rect 1280 1170 1300 1190
rect 1380 1170 1400 1190
rect 1480 1170 1500 1190
rect 1580 1170 1600 1190
rect 1680 1170 1700 1190
rect 1780 1170 1800 1190
rect 1880 1170 1900 1190
rect 1980 1170 2000 1190
rect 30 950 50 970
rect 1080 950 1100 970
rect 2130 950 2150 970
rect 30 820 50 840
rect 1080 820 1100 840
rect 1280 820 1300 840
rect 1380 820 1400 840
rect 1480 820 1500 840
rect 1580 820 1600 840
rect 1680 820 1700 840
rect 1780 820 1800 840
rect 1880 820 1900 840
rect 1980 820 2000 840
rect 2130 820 2150 840
rect 30 -55 50 -35
rect 180 -55 200 -35
rect 280 -55 300 -35
rect 380 -55 400 -35
rect 480 -55 500 -35
rect 580 -55 600 -35
rect 680 -55 700 -35
rect 780 -55 800 -35
rect 880 -55 900 -35
rect 1080 -50 1100 -30
rect 1280 -50 1300 -30
rect 1380 -50 1400 -30
rect 1480 -50 1500 -30
rect 1580 -50 1600 -30
rect 1680 -50 1700 -30
rect 1780 -50 1800 -30
rect 1880 -50 1900 -30
rect 1980 -50 2000 -30
rect 2130 -50 2150 -30
<< locali >>
rect 120 1190 2060 1200
rect 120 1170 180 1190
rect 200 1170 280 1190
rect 300 1170 380 1190
rect 400 1170 480 1190
rect 500 1170 580 1190
rect 600 1170 680 1190
rect 700 1170 780 1190
rect 800 1170 880 1190
rect 900 1170 1280 1190
rect 1300 1170 1380 1190
rect 1400 1170 1480 1190
rect 1500 1170 1580 1190
rect 1600 1170 1680 1190
rect 1700 1170 1780 1190
rect 1800 1170 1880 1190
rect 1900 1170 1980 1190
rect 2000 1170 2060 1190
rect 120 1160 2060 1170
rect -35 1130 60 1140
rect -35 1010 -25 1130
rect 0 1010 30 1130
rect 50 1010 60 1130
rect -35 1000 60 1010
rect 120 1130 160 1160
rect 120 1010 130 1130
rect 150 1010 160 1130
rect 120 1000 160 1010
rect 220 1130 260 1140
rect 220 1010 230 1130
rect 250 1010 260 1130
rect 220 1000 260 1010
rect 320 1130 360 1140
rect 320 1010 330 1130
rect 350 1010 360 1130
rect 320 1000 360 1010
rect 420 1130 460 1140
rect 420 1010 430 1130
rect 450 1010 460 1130
rect 420 1000 460 1010
rect 520 1130 560 1160
rect 520 1010 530 1130
rect 550 1010 560 1130
rect 520 1000 560 1010
rect 620 1130 660 1140
rect 620 1010 630 1130
rect 650 1010 660 1130
rect 620 1000 660 1010
rect 720 1130 760 1140
rect 720 1010 730 1130
rect 750 1010 760 1130
rect 720 1000 760 1010
rect 820 1130 860 1140
rect 820 1010 830 1130
rect 850 1010 860 1130
rect 820 1000 860 1010
rect 920 1130 960 1160
rect 920 1010 930 1130
rect 950 1010 960 1130
rect 920 1000 960 1010
rect 1020 1130 1160 1140
rect 1020 1010 1030 1130
rect 1050 1010 1080 1130
rect 1100 1010 1130 1130
rect 1150 1010 1160 1130
rect 1020 1000 1160 1010
rect 1220 1130 1260 1160
rect 1220 1010 1230 1130
rect 1250 1010 1260 1130
rect 1220 1000 1260 1010
rect 1320 1130 1360 1140
rect 1320 1010 1330 1130
rect 1350 1010 1360 1130
rect 1320 1000 1360 1010
rect 1420 1130 1460 1140
rect 1420 1010 1430 1130
rect 1450 1010 1460 1130
rect 1420 1000 1460 1010
rect 1520 1130 1560 1140
rect 1520 1010 1530 1130
rect 1550 1010 1560 1130
rect 1520 1000 1560 1010
rect 1620 1130 1660 1160
rect 1620 1010 1630 1130
rect 1650 1010 1660 1130
rect 1620 1000 1660 1010
rect 1720 1130 1760 1140
rect 1720 1010 1730 1130
rect 1750 1010 1760 1130
rect 1720 1000 1760 1010
rect 1820 1130 1860 1140
rect 1820 1010 1830 1130
rect 1850 1010 1860 1130
rect 1820 1000 1860 1010
rect 1920 1130 1960 1140
rect 1920 1010 1930 1130
rect 1950 1010 1960 1130
rect 1920 1000 1960 1010
rect 2020 1130 2060 1160
rect 2020 1010 2030 1130
rect 2050 1010 2060 1130
rect 2020 1000 2060 1010
rect 2120 1130 2210 1140
rect 2120 1010 2130 1130
rect 2150 1010 2180 1130
rect 2200 1010 2210 1130
rect 2120 1000 2210 1010
rect 20 970 60 1000
rect 20 950 30 970
rect 50 950 60 970
rect 20 940 60 950
rect 1070 970 1110 1000
rect 1070 950 1080 970
rect 1100 950 1110 970
rect 1070 940 1110 950
rect 2120 970 2160 1000
rect 2120 950 2130 970
rect 2150 950 2160 970
rect 2120 940 2160 950
rect 20 840 60 850
rect 20 820 30 840
rect 50 820 60 840
rect 20 790 60 820
rect 1070 840 1110 850
rect 1070 820 1080 840
rect 1100 820 1110 840
rect 1070 790 1110 820
rect 1220 840 2060 850
rect 1220 820 1280 840
rect 1300 820 1380 840
rect 1400 820 1480 840
rect 1500 820 1580 840
rect 1600 820 1680 840
rect 1700 820 1780 840
rect 1800 820 1880 840
rect 1900 820 1980 840
rect 2000 820 2060 840
rect 1220 810 2060 820
rect -35 780 60 790
rect -35 510 -25 780
rect 0 510 30 780
rect 50 510 60 780
rect -35 500 60 510
rect 120 780 160 790
rect 120 510 130 780
rect 150 510 160 780
rect 120 500 160 510
rect 220 780 260 790
rect 220 510 230 780
rect 250 510 260 780
rect 220 500 260 510
rect 320 780 360 790
rect 320 510 330 780
rect 350 510 360 780
rect 320 500 360 510
rect 420 780 460 790
rect 420 510 430 780
rect 450 510 460 780
rect 420 500 460 510
rect 520 780 560 790
rect 520 510 530 780
rect 550 510 560 780
rect 520 500 560 510
rect 620 780 660 790
rect 620 510 630 780
rect 650 510 660 780
rect 620 500 660 510
rect 720 780 760 790
rect 720 510 730 780
rect 750 510 760 780
rect 720 500 760 510
rect 820 780 860 790
rect 820 510 830 780
rect 850 510 860 780
rect 820 500 860 510
rect 920 780 960 790
rect 920 510 930 780
rect 950 510 960 780
rect 920 500 960 510
rect 1020 780 1160 790
rect 1020 510 1030 780
rect 1050 510 1080 780
rect 1100 510 1130 780
rect 1150 510 1160 780
rect 1020 500 1160 510
rect 1220 780 1260 810
rect 1220 510 1230 780
rect 1250 510 1260 780
rect 1220 500 1260 510
rect 1320 780 1360 790
rect 1320 510 1330 780
rect 1350 510 1360 780
rect 1320 500 1360 510
rect 1420 780 1460 790
rect 1420 510 1430 780
rect 1450 510 1460 780
rect 1420 500 1460 510
rect 1520 780 1560 790
rect 1520 510 1530 780
rect 1550 510 1560 780
rect 1520 500 1560 510
rect 1620 780 1660 810
rect 1620 510 1630 780
rect 1650 510 1660 780
rect 1620 500 1660 510
rect 1720 780 1760 790
rect 1720 510 1730 780
rect 1750 510 1760 780
rect 1720 500 1760 510
rect 1820 780 1860 790
rect 1820 510 1830 780
rect 1850 510 1860 780
rect 1820 500 1860 510
rect 1920 780 1960 790
rect 1920 510 1930 780
rect 1950 510 1960 780
rect 1920 500 1960 510
rect 2020 780 2060 810
rect 2020 510 2030 780
rect 2050 510 2060 780
rect 2020 500 2060 510
rect 2120 840 2160 850
rect 2120 820 2130 840
rect 2150 820 2160 840
rect 2120 790 2160 820
rect 2120 780 2210 790
rect 2120 510 2130 780
rect 2150 510 2180 780
rect 2200 510 2210 780
rect 2120 500 2210 510
rect -35 280 60 290
rect -35 10 -25 280
rect 0 10 30 280
rect 50 10 60 280
rect -35 0 60 10
rect 20 -35 60 0
rect 20 -55 30 -35
rect 50 -55 60 -35
rect 20 -65 60 -55
rect 120 280 160 290
rect 120 10 130 280
rect 150 10 160 280
rect 120 -25 160 10
rect 220 280 260 290
rect 220 10 230 280
rect 250 10 260 280
rect 220 0 260 10
rect 320 280 360 290
rect 320 10 330 280
rect 350 10 360 280
rect 320 0 360 10
rect 420 280 460 290
rect 420 10 430 280
rect 450 10 460 280
rect 420 0 460 10
rect 520 280 560 290
rect 520 10 530 280
rect 550 10 560 280
rect 520 -25 560 10
rect 620 280 660 290
rect 620 10 630 280
rect 650 10 660 280
rect 620 0 660 10
rect 720 280 760 290
rect 720 10 730 280
rect 750 10 760 280
rect 720 0 760 10
rect 820 280 860 290
rect 820 10 830 280
rect 850 10 860 280
rect 820 0 860 10
rect 920 280 960 290
rect 920 10 930 280
rect 950 10 960 280
rect 920 -25 960 10
rect 1020 280 1160 290
rect 1020 10 1030 280
rect 1050 10 1080 280
rect 1100 10 1130 280
rect 1150 10 1160 280
rect 1020 0 1160 10
rect 1220 280 1260 290
rect 1220 10 1230 280
rect 1250 10 1260 280
rect 120 -35 960 -25
rect 120 -55 180 -35
rect 200 -55 280 -35
rect 300 -55 380 -35
rect 400 -55 480 -35
rect 500 -55 580 -35
rect 600 -55 680 -35
rect 700 -55 780 -35
rect 800 -55 880 -35
rect 900 -55 960 -35
rect 120 -65 960 -55
rect 1070 -30 1110 0
rect 1070 -50 1080 -30
rect 1100 -50 1110 -30
rect 1070 -60 1110 -50
rect 1220 -20 1260 10
rect 1320 280 1360 290
rect 1320 10 1330 280
rect 1350 10 1360 280
rect 1320 0 1360 10
rect 1420 280 1460 290
rect 1420 10 1430 280
rect 1450 10 1460 280
rect 1420 0 1460 10
rect 1520 280 1560 290
rect 1520 10 1530 280
rect 1550 10 1560 280
rect 1520 0 1560 10
rect 1620 280 1660 290
rect 1620 10 1630 280
rect 1650 10 1660 280
rect 1620 -20 1660 10
rect 1720 280 1760 290
rect 1720 10 1730 280
rect 1750 10 1760 280
rect 1720 0 1760 10
rect 1820 280 1860 290
rect 1820 10 1830 280
rect 1850 10 1860 280
rect 1820 0 1860 10
rect 1920 280 1960 290
rect 1920 10 1930 280
rect 1950 10 1960 280
rect 1920 0 1960 10
rect 2020 280 2060 290
rect 2020 10 2030 280
rect 2050 10 2060 280
rect 2020 -20 2060 10
rect 1220 -30 2060 -20
rect 1220 -50 1280 -30
rect 1300 -50 1380 -30
rect 1400 -50 1480 -30
rect 1500 -50 1580 -30
rect 1600 -50 1680 -30
rect 1700 -50 1780 -30
rect 1800 -50 1880 -30
rect 1900 -50 1980 -30
rect 2000 -50 2060 -30
rect 1220 -60 2060 -50
rect 2120 280 2210 290
rect 2120 10 2130 280
rect 2150 10 2180 280
rect 2200 10 2210 280
rect 2120 0 2210 10
rect 2120 -30 2160 0
rect 2120 -50 2130 -30
rect 2150 -50 2160 -30
rect 2120 -60 2160 -50
<< viali >>
rect 30 1010 50 1130
rect 230 1010 250 1130
rect 430 1010 450 1130
rect 630 1010 650 1130
rect 830 1010 850 1130
rect 1030 1010 1050 1130
rect 1080 1010 1100 1130
rect 1130 1010 1150 1130
rect 1330 1010 1350 1130
rect 1530 1010 1550 1130
rect 1730 1010 1750 1130
rect 1930 1010 1950 1130
rect 2130 1010 2150 1130
rect 2180 1010 2200 1130
rect -25 510 0 780
rect 1030 510 1050 780
rect 1080 510 1100 780
rect 1130 510 1150 780
rect 1330 510 1350 780
rect 1530 510 1550 780
rect 1730 510 1750 780
rect 1930 510 1950 780
rect 2130 510 2150 780
rect 2180 510 2200 780
rect -25 10 0 280
rect 30 10 50 280
rect 230 10 250 280
rect 430 10 450 280
rect 630 10 650 280
rect 830 10 850 280
rect 1030 10 1050 280
rect 1080 10 1100 280
rect 1130 10 1150 280
rect 1330 10 1350 280
rect 1530 10 1550 280
rect 1730 10 1750 280
rect 1930 10 1950 280
rect 2130 10 2150 280
rect 2180 10 2200 280
<< metal1 >>
rect -60 1130 2235 1140
rect -60 1010 30 1130
rect 50 1010 230 1130
rect 250 1010 430 1130
rect 450 1010 630 1130
rect 650 1010 830 1130
rect 850 1010 1030 1130
rect 1050 1010 1080 1130
rect 1100 1010 1130 1130
rect 1150 1010 1330 1130
rect 1350 1010 1530 1130
rect 1550 1010 1730 1130
rect 1750 1010 1930 1130
rect 1950 1010 2130 1130
rect 2150 1010 2180 1130
rect 2200 1010 2235 1130
rect -60 780 2235 1010
rect -60 510 -25 780
rect 0 510 1030 780
rect 1050 510 1080 780
rect 1100 510 1130 780
rect 1150 510 1330 780
rect 1350 510 1530 780
rect 1550 510 1730 780
rect 1750 510 1930 780
rect 1950 510 2130 780
rect 2150 510 2180 780
rect 2200 510 2235 780
rect -60 505 2235 510
rect -35 280 2210 290
rect -35 10 -25 280
rect 0 10 30 280
rect 50 10 230 280
rect 250 10 430 280
rect 450 10 630 280
rect 650 10 830 280
rect 850 10 1030 280
rect 1050 10 1080 280
rect 1100 10 1130 280
rect 1150 10 1330 280
rect 1350 10 1530 280
rect 1550 10 1730 280
rect 1750 10 1930 280
rect 1950 10 2130 280
rect 2150 10 2180 280
rect 2200 10 2210 280
rect -35 0 2210 10
<< end >>
